LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.SDRNCO_pkg.ALL;

ENTITY SDRNCOLookUpTableGen IS
  PORT( clk                               :   IN    std_logic;
        reset                             :   IN    std_logic;
        enb                               :   IN    std_logic;
        lutaddr                           :   IN    std_logic_vector(17 DOWNTO 0);  -- ufix18
        lutoutput                         :   OUT   std_logic_vector(19 DOWNTO 0)  -- sfix20_En18
        );
END SDRNCOLookUpTableGen;


ARCHITECTURE rtl OF SDRNCOLookUpTableGen IS

  -- Constants
  CONSTANT table_data                     : vector_of_signed20(0 TO 4095) := ( to_signed(16#00000#, 20), to_signed(16#00065#, 20), to_signed(16#000C9#, 20), to_signed(16#0012E#, 20),
                                                                              to_signed(16#00192#, 20), to_signed(16#001F7#, 20), to_signed(16#0025B#, 20), to_signed(16#002C0#, 20),
                                                                              to_signed(16#00324#, 20), to_signed(16#00389#, 20), to_signed(16#003ED#, 20), to_signed(16#00452#, 20),
                                                                              to_signed(16#004B6#, 20), to_signed(16#0051B#, 20), to_signed(16#0057F#, 20), to_signed(16#005E4#, 20),
                                                                              to_signed(16#00648#, 20), to_signed(16#006AD#, 20), to_signed(16#00712#, 20), to_signed(16#00776#, 20),
                                                                              to_signed(16#007DB#, 20), to_signed(16#0083F#, 20), to_signed(16#008A4#, 20), to_signed(16#00908#, 20),
                                                                              to_signed(16#0096D#, 20), to_signed(16#009D1#, 20), to_signed(16#00A36#, 20), to_signed(16#00A9A#, 20),
                                                                              to_signed(16#00AFF#, 20), to_signed(16#00B63#, 20), to_signed(16#00BC8#, 20), to_signed(16#00C2C#, 20),
                                                                              to_signed(16#00C91#, 20), to_signed(16#00CF5#, 20), to_signed(16#00D5A#, 20), to_signed(16#00DBE#, 20),
                                                                              to_signed(16#00E23#, 20), to_signed(16#00E88#, 20), to_signed(16#00EEC#, 20), to_signed(16#00F51#, 20),
                                                                              to_signed(16#00FB5#, 20), to_signed(16#0101A#, 20), to_signed(16#0107E#, 20), to_signed(16#010E3#, 20),
                                                                              to_signed(16#01147#, 20), to_signed(16#011AC#, 20), to_signed(16#01210#, 20), to_signed(16#01275#, 20),
                                                                              to_signed(16#012D9#, 20), to_signed(16#0133E#, 20), to_signed(16#013A2#, 20), to_signed(16#01407#, 20),
                                                                              to_signed(16#0146B#, 20), to_signed(16#014D0#, 20), to_signed(16#01534#, 20), to_signed(16#01599#, 20),
                                                                              to_signed(16#015FD#, 20), to_signed(16#01662#, 20), to_signed(16#016C6#, 20), to_signed(16#0172B#, 20),
                                                                              to_signed(16#0178F#, 20), to_signed(16#017F4#, 20), to_signed(16#01858#, 20), to_signed(16#018BD#, 20),
                                                                              to_signed(16#01921#, 20), to_signed(16#01986#, 20), to_signed(16#019EA#, 20), to_signed(16#01A4F#, 20),
                                                                              to_signed(16#01AB3#, 20), to_signed(16#01B18#, 20), to_signed(16#01B7C#, 20), to_signed(16#01BE1#, 20),
                                                                              to_signed(16#01C45#, 20), to_signed(16#01CAA#, 20), to_signed(16#01D0E#, 20), to_signed(16#01D73#, 20),
                                                                              to_signed(16#01DD7#, 20), to_signed(16#01E3C#, 20), to_signed(16#01EA0#, 20), to_signed(16#01F05#, 20),
                                                                              to_signed(16#01F69#, 20), to_signed(16#01FCE#, 20), to_signed(16#02032#, 20), to_signed(16#02097#, 20),
                                                                              to_signed(16#020FB#, 20), to_signed(16#02160#, 20), to_signed(16#021C4#, 20), to_signed(16#02229#, 20),
                                                                              to_signed(16#0228D#, 20), to_signed(16#022F2#, 20), to_signed(16#02356#, 20), to_signed(16#023BA#, 20),
                                                                              to_signed(16#0241F#, 20), to_signed(16#02483#, 20), to_signed(16#024E8#, 20), to_signed(16#0254C#, 20),
                                                                              to_signed(16#025B1#, 20), to_signed(16#02615#, 20), to_signed(16#0267A#, 20), to_signed(16#026DE#, 20),
                                                                              to_signed(16#02743#, 20), to_signed(16#027A7#, 20), to_signed(16#0280C#, 20), to_signed(16#02870#, 20),
                                                                              to_signed(16#028D4#, 20), to_signed(16#02939#, 20), to_signed(16#0299D#, 20), to_signed(16#02A02#, 20),
                                                                              to_signed(16#02A66#, 20), to_signed(16#02ACB#, 20), to_signed(16#02B2F#, 20), to_signed(16#02B94#, 20),
                                                                              to_signed(16#02BF8#, 20), to_signed(16#02C5C#, 20), to_signed(16#02CC1#, 20), to_signed(16#02D25#, 20),
                                                                              to_signed(16#02D8A#, 20), to_signed(16#02DEE#, 20), to_signed(16#02E53#, 20), to_signed(16#02EB7#, 20),
                                                                              to_signed(16#02F1B#, 20), to_signed(16#02F80#, 20), to_signed(16#02FE4#, 20), to_signed(16#03049#, 20),
                                                                              to_signed(16#030AD#, 20), to_signed(16#03112#, 20), to_signed(16#03176#, 20), to_signed(16#031DA#, 20),
                                                                              to_signed(16#0323F#, 20), to_signed(16#032A3#, 20), to_signed(16#03308#, 20), to_signed(16#0336C#, 20),
                                                                              to_signed(16#033D0#, 20), to_signed(16#03435#, 20), to_signed(16#03499#, 20), to_signed(16#034FE#, 20),
                                                                              to_signed(16#03562#, 20), to_signed(16#035C6#, 20), to_signed(16#0362B#, 20), to_signed(16#0368F#, 20),
                                                                              to_signed(16#036F4#, 20), to_signed(16#03758#, 20), to_signed(16#037BC#, 20), to_signed(16#03821#, 20),
                                                                              to_signed(16#03885#, 20), to_signed(16#038E9#, 20), to_signed(16#0394E#, 20), to_signed(16#039B2#, 20),
                                                                              to_signed(16#03A17#, 20), to_signed(16#03A7B#, 20), to_signed(16#03ADF#, 20), to_signed(16#03B44#, 20),
                                                                              to_signed(16#03BA8#, 20), to_signed(16#03C0C#, 20), to_signed(16#03C71#, 20), to_signed(16#03CD5#, 20),
                                                                              to_signed(16#03D39#, 20), to_signed(16#03D9E#, 20), to_signed(16#03E02#, 20), to_signed(16#03E67#, 20),
                                                                              to_signed(16#03ECB#, 20), to_signed(16#03F2F#, 20), to_signed(16#03F94#, 20), to_signed(16#03FF8#, 20),
                                                                              to_signed(16#0405C#, 20), to_signed(16#040C1#, 20), to_signed(16#04125#, 20), to_signed(16#04189#, 20),
                                                                              to_signed(16#041EE#, 20), to_signed(16#04252#, 20), to_signed(16#042B6#, 20), to_signed(16#0431A#, 20),
                                                                              to_signed(16#0437F#, 20), to_signed(16#043E3#, 20), to_signed(16#04447#, 20), to_signed(16#044AC#, 20),
                                                                              to_signed(16#04510#, 20), to_signed(16#04574#, 20), to_signed(16#045D9#, 20), to_signed(16#0463D#, 20),
                                                                              to_signed(16#046A1#, 20), to_signed(16#04705#, 20), to_signed(16#0476A#, 20), to_signed(16#047CE#, 20),
                                                                              to_signed(16#04832#, 20), to_signed(16#04897#, 20), to_signed(16#048FB#, 20), to_signed(16#0495F#, 20),
                                                                              to_signed(16#049C3#, 20), to_signed(16#04A28#, 20), to_signed(16#04A8C#, 20), to_signed(16#04AF0#, 20),
                                                                              to_signed(16#04B55#, 20), to_signed(16#04BB9#, 20), to_signed(16#04C1D#, 20), to_signed(16#04C81#, 20),
                                                                              to_signed(16#04CE6#, 20), to_signed(16#04D4A#, 20), to_signed(16#04DAE#, 20), to_signed(16#04E12#, 20),
                                                                              to_signed(16#04E76#, 20), to_signed(16#04EDB#, 20), to_signed(16#04F3F#, 20), to_signed(16#04FA3#, 20),
                                                                              to_signed(16#05007#, 20), to_signed(16#0506C#, 20), to_signed(16#050D0#, 20), to_signed(16#05134#, 20),
                                                                              to_signed(16#05198#, 20), to_signed(16#051FC#, 20), to_signed(16#05261#, 20), to_signed(16#052C5#, 20),
                                                                              to_signed(16#05329#, 20), to_signed(16#0538D#, 20), to_signed(16#053F1#, 20), to_signed(16#05456#, 20),
                                                                              to_signed(16#054BA#, 20), to_signed(16#0551E#, 20), to_signed(16#05582#, 20), to_signed(16#055E6#, 20),
                                                                              to_signed(16#0564B#, 20), to_signed(16#056AF#, 20), to_signed(16#05713#, 20), to_signed(16#05777#, 20),
                                                                              to_signed(16#057DB#, 20), to_signed(16#0583F#, 20), to_signed(16#058A4#, 20), to_signed(16#05908#, 20),
                                                                              to_signed(16#0596C#, 20), to_signed(16#059D0#, 20), to_signed(16#05A34#, 20), to_signed(16#05A98#, 20),
                                                                              to_signed(16#05AFC#, 20), to_signed(16#05B61#, 20), to_signed(16#05BC5#, 20), to_signed(16#05C29#, 20),
                                                                              to_signed(16#05C8D#, 20), to_signed(16#05CF1#, 20), to_signed(16#05D55#, 20), to_signed(16#05DB9#, 20),
                                                                              to_signed(16#05E1D#, 20), to_signed(16#05E81#, 20), to_signed(16#05EE6#, 20), to_signed(16#05F4A#, 20),
                                                                              to_signed(16#05FAE#, 20), to_signed(16#06012#, 20), to_signed(16#06076#, 20), to_signed(16#060DA#, 20),
                                                                              to_signed(16#0613E#, 20), to_signed(16#061A2#, 20), to_signed(16#06206#, 20), to_signed(16#0626A#, 20),
                                                                              to_signed(16#062CE#, 20), to_signed(16#06332#, 20), to_signed(16#06397#, 20), to_signed(16#063FB#, 20),
                                                                              to_signed(16#0645F#, 20), to_signed(16#064C3#, 20), to_signed(16#06527#, 20), to_signed(16#0658B#, 20),
                                                                              to_signed(16#065EF#, 20), to_signed(16#06653#, 20), to_signed(16#066B7#, 20), to_signed(16#0671B#, 20),
                                                                              to_signed(16#0677F#, 20), to_signed(16#067E3#, 20), to_signed(16#06847#, 20), to_signed(16#068AB#, 20),
                                                                              to_signed(16#0690F#, 20), to_signed(16#06973#, 20), to_signed(16#069D7#, 20), to_signed(16#06A3B#, 20),
                                                                              to_signed(16#06A9F#, 20), to_signed(16#06B03#, 20), to_signed(16#06B67#, 20), to_signed(16#06BCB#, 20),
                                                                              to_signed(16#06C2F#, 20), to_signed(16#06C93#, 20), to_signed(16#06CF7#, 20), to_signed(16#06D5B#, 20),
                                                                              to_signed(16#06DBF#, 20), to_signed(16#06E23#, 20), to_signed(16#06E87#, 20), to_signed(16#06EEA#, 20),
                                                                              to_signed(16#06F4E#, 20), to_signed(16#06FB2#, 20), to_signed(16#07016#, 20), to_signed(16#0707A#, 20),
                                                                              to_signed(16#070DE#, 20), to_signed(16#07142#, 20), to_signed(16#071A6#, 20), to_signed(16#0720A#, 20),
                                                                              to_signed(16#0726E#, 20), to_signed(16#072D2#, 20), to_signed(16#07336#, 20), to_signed(16#07399#, 20),
                                                                              to_signed(16#073FD#, 20), to_signed(16#07461#, 20), to_signed(16#074C5#, 20), to_signed(16#07529#, 20),
                                                                              to_signed(16#0758D#, 20), to_signed(16#075F1#, 20), to_signed(16#07655#, 20), to_signed(16#076B8#, 20),
                                                                              to_signed(16#0771C#, 20), to_signed(16#07780#, 20), to_signed(16#077E4#, 20), to_signed(16#07848#, 20),
                                                                              to_signed(16#078AC#, 20), to_signed(16#0790F#, 20), to_signed(16#07973#, 20), to_signed(16#079D7#, 20),
                                                                              to_signed(16#07A3B#, 20), to_signed(16#07A9F#, 20), to_signed(16#07B02#, 20), to_signed(16#07B66#, 20),
                                                                              to_signed(16#07BCA#, 20), to_signed(16#07C2E#, 20), to_signed(16#07C92#, 20), to_signed(16#07CF5#, 20),
                                                                              to_signed(16#07D59#, 20), to_signed(16#07DBD#, 20), to_signed(16#07E21#, 20), to_signed(16#07E85#, 20),
                                                                              to_signed(16#07EE8#, 20), to_signed(16#07F4C#, 20), to_signed(16#07FB0#, 20), to_signed(16#08014#, 20),
                                                                              to_signed(16#08077#, 20), to_signed(16#080DB#, 20), to_signed(16#0813F#, 20), to_signed(16#081A2#, 20),
                                                                              to_signed(16#08206#, 20), to_signed(16#0826A#, 20), to_signed(16#082CE#, 20), to_signed(16#08331#, 20),
                                                                              to_signed(16#08395#, 20), to_signed(16#083F9#, 20), to_signed(16#0845C#, 20), to_signed(16#084C0#, 20),
                                                                              to_signed(16#08524#, 20), to_signed(16#08587#, 20), to_signed(16#085EB#, 20), to_signed(16#0864F#, 20),
                                                                              to_signed(16#086B2#, 20), to_signed(16#08716#, 20), to_signed(16#0877A#, 20), to_signed(16#087DD#, 20),
                                                                              to_signed(16#08841#, 20), to_signed(16#088A5#, 20), to_signed(16#08908#, 20), to_signed(16#0896C#, 20),
                                                                              to_signed(16#089D0#, 20), to_signed(16#08A33#, 20), to_signed(16#08A97#, 20), to_signed(16#08AFA#, 20),
                                                                              to_signed(16#08B5E#, 20), to_signed(16#08BC2#, 20), to_signed(16#08C25#, 20), to_signed(16#08C89#, 20),
                                                                              to_signed(16#08CEC#, 20), to_signed(16#08D50#, 20), to_signed(16#08DB3#, 20), to_signed(16#08E17#, 20),
                                                                              to_signed(16#08E7B#, 20), to_signed(16#08EDE#, 20), to_signed(16#08F42#, 20), to_signed(16#08FA5#, 20),
                                                                              to_signed(16#09009#, 20), to_signed(16#0906C#, 20), to_signed(16#090D0#, 20), to_signed(16#09133#, 20),
                                                                              to_signed(16#09197#, 20), to_signed(16#091FA#, 20), to_signed(16#0925E#, 20), to_signed(16#092C1#, 20),
                                                                              to_signed(16#09325#, 20), to_signed(16#09388#, 20), to_signed(16#093EC#, 20), to_signed(16#0944F#, 20),
                                                                              to_signed(16#094B3#, 20), to_signed(16#09516#, 20), to_signed(16#0957A#, 20), to_signed(16#095DD#, 20),
                                                                              to_signed(16#09641#, 20), to_signed(16#096A4#, 20), to_signed(16#09707#, 20), to_signed(16#0976B#, 20),
                                                                              to_signed(16#097CE#, 20), to_signed(16#09832#, 20), to_signed(16#09895#, 20), to_signed(16#098F8#, 20),
                                                                              to_signed(16#0995C#, 20), to_signed(16#099BF#, 20), to_signed(16#09A23#, 20), to_signed(16#09A86#, 20),
                                                                              to_signed(16#09AE9#, 20), to_signed(16#09B4D#, 20), to_signed(16#09BB0#, 20), to_signed(16#09C14#, 20),
                                                                              to_signed(16#09C77#, 20), to_signed(16#09CDA#, 20), to_signed(16#09D3E#, 20), to_signed(16#09DA1#, 20),
                                                                              to_signed(16#09E04#, 20), to_signed(16#09E68#, 20), to_signed(16#09ECB#, 20), to_signed(16#09F2E#, 20),
                                                                              to_signed(16#09F91#, 20), to_signed(16#09FF5#, 20), to_signed(16#0A058#, 20), to_signed(16#0A0BB#, 20),
                                                                              to_signed(16#0A11F#, 20), to_signed(16#0A182#, 20), to_signed(16#0A1E5#, 20), to_signed(16#0A248#, 20),
                                                                              to_signed(16#0A2AC#, 20), to_signed(16#0A30F#, 20), to_signed(16#0A372#, 20), to_signed(16#0A3D5#, 20),
                                                                              to_signed(16#0A439#, 20), to_signed(16#0A49C#, 20), to_signed(16#0A4FF#, 20), to_signed(16#0A562#, 20),
                                                                              to_signed(16#0A5C6#, 20), to_signed(16#0A629#, 20), to_signed(16#0A68C#, 20), to_signed(16#0A6EF#, 20),
                                                                              to_signed(16#0A752#, 20), to_signed(16#0A7B5#, 20), to_signed(16#0A819#, 20), to_signed(16#0A87C#, 20),
                                                                              to_signed(16#0A8DF#, 20), to_signed(16#0A942#, 20), to_signed(16#0A9A5#, 20), to_signed(16#0AA08#, 20),
                                                                              to_signed(16#0AA6C#, 20), to_signed(16#0AACF#, 20), to_signed(16#0AB32#, 20), to_signed(16#0AB95#, 20),
                                                                              to_signed(16#0ABF8#, 20), to_signed(16#0AC5B#, 20), to_signed(16#0ACBE#, 20), to_signed(16#0AD21#, 20),
                                                                              to_signed(16#0AD84#, 20), to_signed(16#0ADE7#, 20), to_signed(16#0AE4B#, 20), to_signed(16#0AEAE#, 20),
                                                                              to_signed(16#0AF11#, 20), to_signed(16#0AF74#, 20), to_signed(16#0AFD7#, 20), to_signed(16#0B03A#, 20),
                                                                              to_signed(16#0B09D#, 20), to_signed(16#0B100#, 20), to_signed(16#0B163#, 20), to_signed(16#0B1C6#, 20),
                                                                              to_signed(16#0B229#, 20), to_signed(16#0B28C#, 20), to_signed(16#0B2EF#, 20), to_signed(16#0B352#, 20),
                                                                              to_signed(16#0B3B5#, 20), to_signed(16#0B418#, 20), to_signed(16#0B47B#, 20), to_signed(16#0B4DE#, 20),
                                                                              to_signed(16#0B541#, 20), to_signed(16#0B5A4#, 20), to_signed(16#0B606#, 20), to_signed(16#0B669#, 20),
                                                                              to_signed(16#0B6CC#, 20), to_signed(16#0B72F#, 20), to_signed(16#0B792#, 20), to_signed(16#0B7F5#, 20),
                                                                              to_signed(16#0B858#, 20), to_signed(16#0B8BB#, 20), to_signed(16#0B91E#, 20), to_signed(16#0B981#, 20),
                                                                              to_signed(16#0B9E3#, 20), to_signed(16#0BA46#, 20), to_signed(16#0BAA9#, 20), to_signed(16#0BB0C#, 20),
                                                                              to_signed(16#0BB6F#, 20), to_signed(16#0BBD2#, 20), to_signed(16#0BC34#, 20), to_signed(16#0BC97#, 20),
                                                                              to_signed(16#0BCFA#, 20), to_signed(16#0BD5D#, 20), to_signed(16#0BDC0#, 20), to_signed(16#0BE22#, 20),
                                                                              to_signed(16#0BE85#, 20), to_signed(16#0BEE8#, 20), to_signed(16#0BF4B#, 20), to_signed(16#0BFAE#, 20),
                                                                              to_signed(16#0C010#, 20), to_signed(16#0C073#, 20), to_signed(16#0C0D6#, 20), to_signed(16#0C138#, 20),
                                                                              to_signed(16#0C19B#, 20), to_signed(16#0C1FE#, 20), to_signed(16#0C261#, 20), to_signed(16#0C2C3#, 20),
                                                                              to_signed(16#0C326#, 20), to_signed(16#0C389#, 20), to_signed(16#0C3EB#, 20), to_signed(16#0C44E#, 20),
                                                                              to_signed(16#0C4B1#, 20), to_signed(16#0C513#, 20), to_signed(16#0C576#, 20), to_signed(16#0C5D9#, 20),
                                                                              to_signed(16#0C63B#, 20), to_signed(16#0C69E#, 20), to_signed(16#0C701#, 20), to_signed(16#0C763#, 20),
                                                                              to_signed(16#0C7C6#, 20), to_signed(16#0C828#, 20), to_signed(16#0C88B#, 20), to_signed(16#0C8EE#, 20),
                                                                              to_signed(16#0C950#, 20), to_signed(16#0C9B3#, 20), to_signed(16#0CA15#, 20), to_signed(16#0CA78#, 20),
                                                                              to_signed(16#0CADA#, 20), to_signed(16#0CB3D#, 20), to_signed(16#0CB9F#, 20), to_signed(16#0CC02#, 20),
                                                                              to_signed(16#0CC64#, 20), to_signed(16#0CCC7#, 20), to_signed(16#0CD29#, 20), to_signed(16#0CD8C#, 20),
                                                                              to_signed(16#0CDEE#, 20), to_signed(16#0CE51#, 20), to_signed(16#0CEB3#, 20), to_signed(16#0CF16#, 20),
                                                                              to_signed(16#0CF78#, 20), to_signed(16#0CFDB#, 20), to_signed(16#0D03D#, 20), to_signed(16#0D0A0#, 20),
                                                                              to_signed(16#0D102#, 20), to_signed(16#0D164#, 20), to_signed(16#0D1C7#, 20), to_signed(16#0D229#, 20),
                                                                              to_signed(16#0D28C#, 20), to_signed(16#0D2EE#, 20), to_signed(16#0D350#, 20), to_signed(16#0D3B3#, 20),
                                                                              to_signed(16#0D415#, 20), to_signed(16#0D477#, 20), to_signed(16#0D4DA#, 20), to_signed(16#0D53C#, 20),
                                                                              to_signed(16#0D59E#, 20), to_signed(16#0D601#, 20), to_signed(16#0D663#, 20), to_signed(16#0D6C5#, 20),
                                                                              to_signed(16#0D728#, 20), to_signed(16#0D78A#, 20), to_signed(16#0D7EC#, 20), to_signed(16#0D84E#, 20),
                                                                              to_signed(16#0D8B1#, 20), to_signed(16#0D913#, 20), to_signed(16#0D975#, 20), to_signed(16#0D9D7#, 20),
                                                                              to_signed(16#0DA3A#, 20), to_signed(16#0DA9C#, 20), to_signed(16#0DAFE#, 20), to_signed(16#0DB60#, 20),
                                                                              to_signed(16#0DBC2#, 20), to_signed(16#0DC25#, 20), to_signed(16#0DC87#, 20), to_signed(16#0DCE9#, 20),
                                                                              to_signed(16#0DD4B#, 20), to_signed(16#0DDAD#, 20), to_signed(16#0DE0F#, 20), to_signed(16#0DE72#, 20),
                                                                              to_signed(16#0DED4#, 20), to_signed(16#0DF36#, 20), to_signed(16#0DF98#, 20), to_signed(16#0DFFA#, 20),
                                                                              to_signed(16#0E05C#, 20), to_signed(16#0E0BE#, 20), to_signed(16#0E120#, 20), to_signed(16#0E182#, 20),
                                                                              to_signed(16#0E1E4#, 20), to_signed(16#0E246#, 20), to_signed(16#0E2A8#, 20), to_signed(16#0E30A#, 20),
                                                                              to_signed(16#0E36D#, 20), to_signed(16#0E3CF#, 20), to_signed(16#0E431#, 20), to_signed(16#0E493#, 20),
                                                                              to_signed(16#0E4F5#, 20), to_signed(16#0E557#, 20), to_signed(16#0E5B8#, 20), to_signed(16#0E61A#, 20),
                                                                              to_signed(16#0E67C#, 20), to_signed(16#0E6DE#, 20), to_signed(16#0E740#, 20), to_signed(16#0E7A2#, 20),
                                                                              to_signed(16#0E804#, 20), to_signed(16#0E866#, 20), to_signed(16#0E8C8#, 20), to_signed(16#0E92A#, 20),
                                                                              to_signed(16#0E98C#, 20), to_signed(16#0E9EE#, 20), to_signed(16#0EA4F#, 20), to_signed(16#0EAB1#, 20),
                                                                              to_signed(16#0EB13#, 20), to_signed(16#0EB75#, 20), to_signed(16#0EBD7#, 20), to_signed(16#0EC39#, 20),
                                                                              to_signed(16#0EC9A#, 20), to_signed(16#0ECFC#, 20), to_signed(16#0ED5E#, 20), to_signed(16#0EDC0#, 20),
                                                                              to_signed(16#0EE22#, 20), to_signed(16#0EE83#, 20), to_signed(16#0EEE5#, 20), to_signed(16#0EF47#, 20),
                                                                              to_signed(16#0EFA9#, 20), to_signed(16#0F00A#, 20), to_signed(16#0F06C#, 20), to_signed(16#0F0CE#, 20),
                                                                              to_signed(16#0F130#, 20), to_signed(16#0F191#, 20), to_signed(16#0F1F3#, 20), to_signed(16#0F255#, 20),
                                                                              to_signed(16#0F2B6#, 20), to_signed(16#0F318#, 20), to_signed(16#0F37A#, 20), to_signed(16#0F3DB#, 20),
                                                                              to_signed(16#0F43D#, 20), to_signed(16#0F49F#, 20), to_signed(16#0F500#, 20), to_signed(16#0F562#, 20),
                                                                              to_signed(16#0F5C3#, 20), to_signed(16#0F625#, 20), to_signed(16#0F687#, 20), to_signed(16#0F6E8#, 20),
                                                                              to_signed(16#0F74A#, 20), to_signed(16#0F7AB#, 20), to_signed(16#0F80D#, 20), to_signed(16#0F86E#, 20),
                                                                              to_signed(16#0F8D0#, 20), to_signed(16#0F931#, 20), to_signed(16#0F993#, 20), to_signed(16#0F9F4#, 20),
                                                                              to_signed(16#0FA56#, 20), to_signed(16#0FAB7#, 20), to_signed(16#0FB19#, 20), to_signed(16#0FB7A#, 20),
                                                                              to_signed(16#0FBDC#, 20), to_signed(16#0FC3D#, 20), to_signed(16#0FC9F#, 20), to_signed(16#0FD00#, 20),
                                                                              to_signed(16#0FD61#, 20), to_signed(16#0FDC3#, 20), to_signed(16#0FE24#, 20), to_signed(16#0FE86#, 20),
                                                                              to_signed(16#0FEE7#, 20), to_signed(16#0FF48#, 20), to_signed(16#0FFAA#, 20), to_signed(16#1000B#, 20),
                                                                              to_signed(16#1006C#, 20), to_signed(16#100CE#, 20), to_signed(16#1012F#, 20), to_signed(16#10190#, 20),
                                                                              to_signed(16#101F2#, 20), to_signed(16#10253#, 20), to_signed(16#102B4#, 20), to_signed(16#10315#, 20),
                                                                              to_signed(16#10377#, 20), to_signed(16#103D8#, 20), to_signed(16#10439#, 20), to_signed(16#1049A#, 20),
                                                                              to_signed(16#104FC#, 20), to_signed(16#1055D#, 20), to_signed(16#105BE#, 20), to_signed(16#1061F#, 20),
                                                                              to_signed(16#10680#, 20), to_signed(16#106E1#, 20), to_signed(16#10743#, 20), to_signed(16#107A4#, 20),
                                                                              to_signed(16#10805#, 20), to_signed(16#10866#, 20), to_signed(16#108C7#, 20), to_signed(16#10928#, 20),
                                                                              to_signed(16#10989#, 20), to_signed(16#109EA#, 20), to_signed(16#10A4B#, 20), to_signed(16#10AAD#, 20),
                                                                              to_signed(16#10B0E#, 20), to_signed(16#10B6F#, 20), to_signed(16#10BD0#, 20), to_signed(16#10C31#, 20),
                                                                              to_signed(16#10C92#, 20), to_signed(16#10CF3#, 20), to_signed(16#10D54#, 20), to_signed(16#10DB5#, 20),
                                                                              to_signed(16#10E16#, 20), to_signed(16#10E77#, 20), to_signed(16#10ED8#, 20), to_signed(16#10F39#, 20),
                                                                              to_signed(16#10F9A#, 20), to_signed(16#10FFA#, 20), to_signed(16#1105B#, 20), to_signed(16#110BC#, 20),
                                                                              to_signed(16#1111D#, 20), to_signed(16#1117E#, 20), to_signed(16#111DF#, 20), to_signed(16#11240#, 20),
                                                                              to_signed(16#112A1#, 20), to_signed(16#11301#, 20), to_signed(16#11362#, 20), to_signed(16#113C3#, 20),
                                                                              to_signed(16#11424#, 20), to_signed(16#11485#, 20), to_signed(16#114E6#, 20), to_signed(16#11546#, 20),
                                                                              to_signed(16#115A7#, 20), to_signed(16#11608#, 20), to_signed(16#11669#, 20), to_signed(16#116C9#, 20),
                                                                              to_signed(16#1172A#, 20), to_signed(16#1178B#, 20), to_signed(16#117EB#, 20), to_signed(16#1184C#, 20),
                                                                              to_signed(16#118AD#, 20), to_signed(16#1190E#, 20), to_signed(16#1196E#, 20), to_signed(16#119CF#, 20),
                                                                              to_signed(16#11A2F#, 20), to_signed(16#11A90#, 20), to_signed(16#11AF1#, 20), to_signed(16#11B51#, 20),
                                                                              to_signed(16#11BB2#, 20), to_signed(16#11C13#, 20), to_signed(16#11C73#, 20), to_signed(16#11CD4#, 20),
                                                                              to_signed(16#11D34#, 20), to_signed(16#11D95#, 20), to_signed(16#11DF5#, 20), to_signed(16#11E56#, 20),
                                                                              to_signed(16#11EB6#, 20), to_signed(16#11F17#, 20), to_signed(16#11F77#, 20), to_signed(16#11FD8#, 20),
                                                                              to_signed(16#12038#, 20), to_signed(16#12099#, 20), to_signed(16#120F9#, 20), to_signed(16#1215A#, 20),
                                                                              to_signed(16#121BA#, 20), to_signed(16#1221B#, 20), to_signed(16#1227B#, 20), to_signed(16#122DB#, 20),
                                                                              to_signed(16#1233C#, 20), to_signed(16#1239C#, 20), to_signed(16#123FC#, 20), to_signed(16#1245D#, 20),
                                                                              to_signed(16#124BD#, 20), to_signed(16#1251D#, 20), to_signed(16#1257E#, 20), to_signed(16#125DE#, 20),
                                                                              to_signed(16#1263E#, 20), to_signed(16#1269F#, 20), to_signed(16#126FF#, 20), to_signed(16#1275F#, 20),
                                                                              to_signed(16#127BF#, 20), to_signed(16#12820#, 20), to_signed(16#12880#, 20), to_signed(16#128E0#, 20),
                                                                              to_signed(16#12940#, 20), to_signed(16#129A1#, 20), to_signed(16#12A01#, 20), to_signed(16#12A61#, 20),
                                                                              to_signed(16#12AC1#, 20), to_signed(16#12B21#, 20), to_signed(16#12B81#, 20), to_signed(16#12BE2#, 20),
                                                                              to_signed(16#12C42#, 20), to_signed(16#12CA2#, 20), to_signed(16#12D02#, 20), to_signed(16#12D62#, 20),
                                                                              to_signed(16#12DC2#, 20), to_signed(16#12E22#, 20), to_signed(16#12E82#, 20), to_signed(16#12EE2#, 20),
                                                                              to_signed(16#12F42#, 20), to_signed(16#12FA2#, 20), to_signed(16#13002#, 20), to_signed(16#13062#, 20),
                                                                              to_signed(16#130C2#, 20), to_signed(16#13122#, 20), to_signed(16#13182#, 20), to_signed(16#131E2#, 20),
                                                                              to_signed(16#13242#, 20), to_signed(16#132A2#, 20), to_signed(16#13302#, 20), to_signed(16#13362#, 20),
                                                                              to_signed(16#133C2#, 20), to_signed(16#13421#, 20), to_signed(16#13481#, 20), to_signed(16#134E1#, 20),
                                                                              to_signed(16#13541#, 20), to_signed(16#135A1#, 20), to_signed(16#13601#, 20), to_signed(16#13661#, 20),
                                                                              to_signed(16#136C0#, 20), to_signed(16#13720#, 20), to_signed(16#13780#, 20), to_signed(16#137E0#, 20),
                                                                              to_signed(16#1383F#, 20), to_signed(16#1389F#, 20), to_signed(16#138FF#, 20), to_signed(16#1395F#, 20),
                                                                              to_signed(16#139BE#, 20), to_signed(16#13A1E#, 20), to_signed(16#13A7E#, 20), to_signed(16#13ADD#, 20),
                                                                              to_signed(16#13B3D#, 20), to_signed(16#13B9D#, 20), to_signed(16#13BFC#, 20), to_signed(16#13C5C#, 20),
                                                                              to_signed(16#13CBB#, 20), to_signed(16#13D1B#, 20), to_signed(16#13D7B#, 20), to_signed(16#13DDA#, 20),
                                                                              to_signed(16#13E3A#, 20), to_signed(16#13E99#, 20), to_signed(16#13EF9#, 20), to_signed(16#13F58#, 20),
                                                                              to_signed(16#13FB8#, 20), to_signed(16#14017#, 20), to_signed(16#14077#, 20), to_signed(16#140D6#, 20),
                                                                              to_signed(16#14136#, 20), to_signed(16#14195#, 20), to_signed(16#141F5#, 20), to_signed(16#14254#, 20),
                                                                              to_signed(16#142B4#, 20), to_signed(16#14313#, 20), to_signed(16#14372#, 20), to_signed(16#143D2#, 20),
                                                                              to_signed(16#14431#, 20), to_signed(16#14490#, 20), to_signed(16#144F0#, 20), to_signed(16#1454F#, 20),
                                                                              to_signed(16#145AE#, 20), to_signed(16#1460E#, 20), to_signed(16#1466D#, 20), to_signed(16#146CC#, 20),
                                                                              to_signed(16#1472C#, 20), to_signed(16#1478B#, 20), to_signed(16#147EA#, 20), to_signed(16#14849#, 20),
                                                                              to_signed(16#148A8#, 20), to_signed(16#14908#, 20), to_signed(16#14967#, 20), to_signed(16#149C6#, 20),
                                                                              to_signed(16#14A25#, 20), to_signed(16#14A84#, 20), to_signed(16#14AE4#, 20), to_signed(16#14B43#, 20),
                                                                              to_signed(16#14BA2#, 20), to_signed(16#14C01#, 20), to_signed(16#14C60#, 20), to_signed(16#14CBF#, 20),
                                                                              to_signed(16#14D1E#, 20), to_signed(16#14D7D#, 20), to_signed(16#14DDC#, 20), to_signed(16#14E3B#, 20),
                                                                              to_signed(16#14E9A#, 20), to_signed(16#14EF9#, 20), to_signed(16#14F58#, 20), to_signed(16#14FB7#, 20),
                                                                              to_signed(16#15016#, 20), to_signed(16#15075#, 20), to_signed(16#150D4#, 20), to_signed(16#15133#, 20),
                                                                              to_signed(16#15192#, 20), to_signed(16#151F1#, 20), to_signed(16#15250#, 20), to_signed(16#152AF#, 20),
                                                                              to_signed(16#1530E#, 20), to_signed(16#1536C#, 20), to_signed(16#153CB#, 20), to_signed(16#1542A#, 20),
                                                                              to_signed(16#15489#, 20), to_signed(16#154E8#, 20), to_signed(16#15546#, 20), to_signed(16#155A5#, 20),
                                                                              to_signed(16#15604#, 20), to_signed(16#15663#, 20), to_signed(16#156C1#, 20), to_signed(16#15720#, 20),
                                                                              to_signed(16#1577F#, 20), to_signed(16#157DE#, 20), to_signed(16#1583C#, 20), to_signed(16#1589B#, 20),
                                                                              to_signed(16#158FA#, 20), to_signed(16#15958#, 20), to_signed(16#159B7#, 20), to_signed(16#15A16#, 20),
                                                                              to_signed(16#15A74#, 20), to_signed(16#15AD3#, 20), to_signed(16#15B31#, 20), to_signed(16#15B90#, 20),
                                                                              to_signed(16#15BEE#, 20), to_signed(16#15C4D#, 20), to_signed(16#15CAC#, 20), to_signed(16#15D0A#, 20),
                                                                              to_signed(16#15D69#, 20), to_signed(16#15DC7#, 20), to_signed(16#15E26#, 20), to_signed(16#15E84#, 20),
                                                                              to_signed(16#15EE2#, 20), to_signed(16#15F41#, 20), to_signed(16#15F9F#, 20), to_signed(16#15FFE#, 20),
                                                                              to_signed(16#1605C#, 20), to_signed(16#160BB#, 20), to_signed(16#16119#, 20), to_signed(16#16177#, 20),
                                                                              to_signed(16#161D6#, 20), to_signed(16#16234#, 20), to_signed(16#16292#, 20), to_signed(16#162F1#, 20),
                                                                              to_signed(16#1634F#, 20), to_signed(16#163AD#, 20), to_signed(16#1640B#, 20), to_signed(16#1646A#, 20),
                                                                              to_signed(16#164C8#, 20), to_signed(16#16526#, 20), to_signed(16#16584#, 20), to_signed(16#165E3#, 20),
                                                                              to_signed(16#16641#, 20), to_signed(16#1669F#, 20), to_signed(16#166FD#, 20), to_signed(16#1675B#, 20),
                                                                              to_signed(16#167B9#, 20), to_signed(16#16817#, 20), to_signed(16#16876#, 20), to_signed(16#168D4#, 20),
                                                                              to_signed(16#16932#, 20), to_signed(16#16990#, 20), to_signed(16#169EE#, 20), to_signed(16#16A4C#, 20),
                                                                              to_signed(16#16AAA#, 20), to_signed(16#16B08#, 20), to_signed(16#16B66#, 20), to_signed(16#16BC4#, 20),
                                                                              to_signed(16#16C22#, 20), to_signed(16#16C80#, 20), to_signed(16#16CDE#, 20), to_signed(16#16D3C#, 20),
                                                                              to_signed(16#16D9A#, 20), to_signed(16#16DF7#, 20), to_signed(16#16E55#, 20), to_signed(16#16EB3#, 20),
                                                                              to_signed(16#16F11#, 20), to_signed(16#16F6F#, 20), to_signed(16#16FCD#, 20), to_signed(16#1702B#, 20),
                                                                              to_signed(16#17088#, 20), to_signed(16#170E6#, 20), to_signed(16#17144#, 20), to_signed(16#171A2#, 20),
                                                                              to_signed(16#171FF#, 20), to_signed(16#1725D#, 20), to_signed(16#172BB#, 20), to_signed(16#17319#, 20),
                                                                              to_signed(16#17376#, 20), to_signed(16#173D4#, 20), to_signed(16#17432#, 20), to_signed(16#1748F#, 20),
                                                                              to_signed(16#174ED#, 20), to_signed(16#1754A#, 20), to_signed(16#175A8#, 20), to_signed(16#17606#, 20),
                                                                              to_signed(16#17663#, 20), to_signed(16#176C1#, 20), to_signed(16#1771E#, 20), to_signed(16#1777C#, 20),
                                                                              to_signed(16#177D9#, 20), to_signed(16#17837#, 20), to_signed(16#17894#, 20), to_signed(16#178F2#, 20),
                                                                              to_signed(16#1794F#, 20), to_signed(16#179AD#, 20), to_signed(16#17A0A#, 20), to_signed(16#17A68#, 20),
                                                                              to_signed(16#17AC5#, 20), to_signed(16#17B22#, 20), to_signed(16#17B80#, 20), to_signed(16#17BDD#, 20),
                                                                              to_signed(16#17C3B#, 20), to_signed(16#17C98#, 20), to_signed(16#17CF5#, 20), to_signed(16#17D53#, 20),
                                                                              to_signed(16#17DB0#, 20), to_signed(16#17E0D#, 20), to_signed(16#17E6A#, 20), to_signed(16#17EC8#, 20),
                                                                              to_signed(16#17F25#, 20), to_signed(16#17F82#, 20), to_signed(16#17FDF#, 20), to_signed(16#1803C#, 20),
                                                                              to_signed(16#1809A#, 20), to_signed(16#180F7#, 20), to_signed(16#18154#, 20), to_signed(16#181B1#, 20),
                                                                              to_signed(16#1820E#, 20), to_signed(16#1826B#, 20), to_signed(16#182C8#, 20), to_signed(16#18326#, 20),
                                                                              to_signed(16#18383#, 20), to_signed(16#183E0#, 20), to_signed(16#1843D#, 20), to_signed(16#1849A#, 20),
                                                                              to_signed(16#184F7#, 20), to_signed(16#18554#, 20), to_signed(16#185B1#, 20), to_signed(16#1860E#, 20),
                                                                              to_signed(16#1866B#, 20), to_signed(16#186C7#, 20), to_signed(16#18724#, 20), to_signed(16#18781#, 20),
                                                                              to_signed(16#187DE#, 20), to_signed(16#1883B#, 20), to_signed(16#18898#, 20), to_signed(16#188F5#, 20),
                                                                              to_signed(16#18952#, 20), to_signed(16#189AE#, 20), to_signed(16#18A0B#, 20), to_signed(16#18A68#, 20),
                                                                              to_signed(16#18AC5#, 20), to_signed(16#18B21#, 20), to_signed(16#18B7E#, 20), to_signed(16#18BDB#, 20),
                                                                              to_signed(16#18C38#, 20), to_signed(16#18C94#, 20), to_signed(16#18CF1#, 20), to_signed(16#18D4E#, 20),
                                                                              to_signed(16#18DAA#, 20), to_signed(16#18E07#, 20), to_signed(16#18E64#, 20), to_signed(16#18EC0#, 20),
                                                                              to_signed(16#18F1D#, 20), to_signed(16#18F79#, 20), to_signed(16#18FD6#, 20), to_signed(16#19032#, 20),
                                                                              to_signed(16#1908F#, 20), to_signed(16#190EB#, 20), to_signed(16#19148#, 20), to_signed(16#191A4#, 20),
                                                                              to_signed(16#19201#, 20), to_signed(16#1925D#, 20), to_signed(16#192BA#, 20), to_signed(16#19316#, 20),
                                                                              to_signed(16#19373#, 20), to_signed(16#193CF#, 20), to_signed(16#1942B#, 20), to_signed(16#19488#, 20),
                                                                              to_signed(16#194E4#, 20), to_signed(16#19540#, 20), to_signed(16#1959D#, 20), to_signed(16#195F9#, 20),
                                                                              to_signed(16#19655#, 20), to_signed(16#196B2#, 20), to_signed(16#1970E#, 20), to_signed(16#1976A#, 20),
                                                                              to_signed(16#197C6#, 20), to_signed(16#19823#, 20), to_signed(16#1987F#, 20), to_signed(16#198DB#, 20),
                                                                              to_signed(16#19937#, 20), to_signed(16#19993#, 20), to_signed(16#199EF#, 20), to_signed(16#19A4B#, 20),
                                                                              to_signed(16#19AA8#, 20), to_signed(16#19B04#, 20), to_signed(16#19B60#, 20), to_signed(16#19BBC#, 20),
                                                                              to_signed(16#19C18#, 20), to_signed(16#19C74#, 20), to_signed(16#19CD0#, 20), to_signed(16#19D2C#, 20),
                                                                              to_signed(16#19D88#, 20), to_signed(16#19DE4#, 20), to_signed(16#19E40#, 20), to_signed(16#19E9C#, 20),
                                                                              to_signed(16#19EF8#, 20), to_signed(16#19F53#, 20), to_signed(16#19FAF#, 20), to_signed(16#1A00B#, 20),
                                                                              to_signed(16#1A067#, 20), to_signed(16#1A0C3#, 20), to_signed(16#1A11F#, 20), to_signed(16#1A17B#, 20),
                                                                              to_signed(16#1A1D6#, 20), to_signed(16#1A232#, 20), to_signed(16#1A28E#, 20), to_signed(16#1A2EA#, 20),
                                                                              to_signed(16#1A345#, 20), to_signed(16#1A3A1#, 20), to_signed(16#1A3FD#, 20), to_signed(16#1A458#, 20),
                                                                              to_signed(16#1A4B4#, 20), to_signed(16#1A510#, 20), to_signed(16#1A56B#, 20), to_signed(16#1A5C7#, 20),
                                                                              to_signed(16#1A623#, 20), to_signed(16#1A67E#, 20), to_signed(16#1A6DA#, 20), to_signed(16#1A735#, 20),
                                                                              to_signed(16#1A791#, 20), to_signed(16#1A7EC#, 20), to_signed(16#1A848#, 20), to_signed(16#1A8A3#, 20),
                                                                              to_signed(16#1A8FF#, 20), to_signed(16#1A95A#, 20), to_signed(16#1A9B6#, 20), to_signed(16#1AA11#, 20),
                                                                              to_signed(16#1AA6D#, 20), to_signed(16#1AAC8#, 20), to_signed(16#1AB23#, 20), to_signed(16#1AB7F#, 20),
                                                                              to_signed(16#1ABDA#, 20), to_signed(16#1AC35#, 20), to_signed(16#1AC91#, 20), to_signed(16#1ACEC#, 20),
                                                                              to_signed(16#1AD47#, 20), to_signed(16#1ADA2#, 20), to_signed(16#1ADFE#, 20), to_signed(16#1AE59#, 20),
                                                                              to_signed(16#1AEB4#, 20), to_signed(16#1AF0F#, 20), to_signed(16#1AF6B#, 20), to_signed(16#1AFC6#, 20),
                                                                              to_signed(16#1B021#, 20), to_signed(16#1B07C#, 20), to_signed(16#1B0D7#, 20), to_signed(16#1B132#, 20),
                                                                              to_signed(16#1B18D#, 20), to_signed(16#1B1E8#, 20), to_signed(16#1B243#, 20), to_signed(16#1B29E#, 20),
                                                                              to_signed(16#1B2F9#, 20), to_signed(16#1B354#, 20), to_signed(16#1B3AF#, 20), to_signed(16#1B40A#, 20),
                                                                              to_signed(16#1B465#, 20), to_signed(16#1B4C0#, 20), to_signed(16#1B51B#, 20), to_signed(16#1B576#, 20),
                                                                              to_signed(16#1B5D1#, 20), to_signed(16#1B62C#, 20), to_signed(16#1B687#, 20), to_signed(16#1B6E2#, 20),
                                                                              to_signed(16#1B73C#, 20), to_signed(16#1B797#, 20), to_signed(16#1B7F2#, 20), to_signed(16#1B84D#, 20),
                                                                              to_signed(16#1B8A8#, 20), to_signed(16#1B902#, 20), to_signed(16#1B95D#, 20), to_signed(16#1B9B8#, 20),
                                                                              to_signed(16#1BA12#, 20), to_signed(16#1BA6D#, 20), to_signed(16#1BAC8#, 20), to_signed(16#1BB22#, 20),
                                                                              to_signed(16#1BB7D#, 20), to_signed(16#1BBD8#, 20), to_signed(16#1BC32#, 20), to_signed(16#1BC8D#, 20),
                                                                              to_signed(16#1BCE7#, 20), to_signed(16#1BD42#, 20), to_signed(16#1BD9C#, 20), to_signed(16#1BDF7#, 20),
                                                                              to_signed(16#1BE51#, 20), to_signed(16#1BEAC#, 20), to_signed(16#1BF06#, 20), to_signed(16#1BF61#, 20),
                                                                              to_signed(16#1BFBB#, 20), to_signed(16#1C016#, 20), to_signed(16#1C070#, 20), to_signed(16#1C0CA#, 20),
                                                                              to_signed(16#1C125#, 20), to_signed(16#1C17F#, 20), to_signed(16#1C1D9#, 20), to_signed(16#1C234#, 20),
                                                                              to_signed(16#1C28E#, 20), to_signed(16#1C2E8#, 20), to_signed(16#1C342#, 20), to_signed(16#1C39D#, 20),
                                                                              to_signed(16#1C3F7#, 20), to_signed(16#1C451#, 20), to_signed(16#1C4AB#, 20), to_signed(16#1C505#, 20),
                                                                              to_signed(16#1C560#, 20), to_signed(16#1C5BA#, 20), to_signed(16#1C614#, 20), to_signed(16#1C66E#, 20),
                                                                              to_signed(16#1C6C8#, 20), to_signed(16#1C722#, 20), to_signed(16#1C77C#, 20), to_signed(16#1C7D6#, 20),
                                                                              to_signed(16#1C830#, 20), to_signed(16#1C88A#, 20), to_signed(16#1C8E4#, 20), to_signed(16#1C93E#, 20),
                                                                              to_signed(16#1C998#, 20), to_signed(16#1C9F2#, 20), to_signed(16#1CA4C#, 20), to_signed(16#1CAA6#, 20),
                                                                              to_signed(16#1CB00#, 20), to_signed(16#1CB59#, 20), to_signed(16#1CBB3#, 20), to_signed(16#1CC0D#, 20),
                                                                              to_signed(16#1CC67#, 20), to_signed(16#1CCC1#, 20), to_signed(16#1CD1A#, 20), to_signed(16#1CD74#, 20),
                                                                              to_signed(16#1CDCE#, 20), to_signed(16#1CE28#, 20), to_signed(16#1CE81#, 20), to_signed(16#1CEDB#, 20),
                                                                              to_signed(16#1CF35#, 20), to_signed(16#1CF8E#, 20), to_signed(16#1CFE8#, 20), to_signed(16#1D042#, 20),
                                                                              to_signed(16#1D09B#, 20), to_signed(16#1D0F5#, 20), to_signed(16#1D14E#, 20), to_signed(16#1D1A8#, 20),
                                                                              to_signed(16#1D201#, 20), to_signed(16#1D25B#, 20), to_signed(16#1D2B4#, 20), to_signed(16#1D30E#, 20),
                                                                              to_signed(16#1D367#, 20), to_signed(16#1D3C1#, 20), to_signed(16#1D41A#, 20), to_signed(16#1D474#, 20),
                                                                              to_signed(16#1D4CD#, 20), to_signed(16#1D526#, 20), to_signed(16#1D580#, 20), to_signed(16#1D5D9#, 20),
                                                                              to_signed(16#1D632#, 20), to_signed(16#1D68C#, 20), to_signed(16#1D6E5#, 20), to_signed(16#1D73E#, 20),
                                                                              to_signed(16#1D797#, 20), to_signed(16#1D7F1#, 20), to_signed(16#1D84A#, 20), to_signed(16#1D8A3#, 20),
                                                                              to_signed(16#1D8FC#, 20), to_signed(16#1D955#, 20), to_signed(16#1D9AF#, 20), to_signed(16#1DA08#, 20),
                                                                              to_signed(16#1DA61#, 20), to_signed(16#1DABA#, 20), to_signed(16#1DB13#, 20), to_signed(16#1DB6C#, 20),
                                                                              to_signed(16#1DBC5#, 20), to_signed(16#1DC1E#, 20), to_signed(16#1DC77#, 20), to_signed(16#1DCD0#, 20),
                                                                              to_signed(16#1DD29#, 20), to_signed(16#1DD82#, 20), to_signed(16#1DDDB#, 20), to_signed(16#1DE34#, 20),
                                                                              to_signed(16#1DE8D#, 20), to_signed(16#1DEE5#, 20), to_signed(16#1DF3E#, 20), to_signed(16#1DF97#, 20),
                                                                              to_signed(16#1DFF0#, 20), to_signed(16#1E049#, 20), to_signed(16#1E0A2#, 20), to_signed(16#1E0FA#, 20),
                                                                              to_signed(16#1E153#, 20), to_signed(16#1E1AC#, 20), to_signed(16#1E204#, 20), to_signed(16#1E25D#, 20),
                                                                              to_signed(16#1E2B6#, 20), to_signed(16#1E30E#, 20), to_signed(16#1E367#, 20), to_signed(16#1E3C0#, 20),
                                                                              to_signed(16#1E418#, 20), to_signed(16#1E471#, 20), to_signed(16#1E4C9#, 20), to_signed(16#1E522#, 20),
                                                                              to_signed(16#1E57B#, 20), to_signed(16#1E5D3#, 20), to_signed(16#1E62C#, 20), to_signed(16#1E684#, 20),
                                                                              to_signed(16#1E6DC#, 20), to_signed(16#1E735#, 20), to_signed(16#1E78D#, 20), to_signed(16#1E7E6#, 20),
                                                                              to_signed(16#1E83E#, 20), to_signed(16#1E896#, 20), to_signed(16#1E8EF#, 20), to_signed(16#1E947#, 20),
                                                                              to_signed(16#1E99F#, 20), to_signed(16#1E9F8#, 20), to_signed(16#1EA50#, 20), to_signed(16#1EAA8#, 20),
                                                                              to_signed(16#1EB00#, 20), to_signed(16#1EB59#, 20), to_signed(16#1EBB1#, 20), to_signed(16#1EC09#, 20),
                                                                              to_signed(16#1EC61#, 20), to_signed(16#1ECB9#, 20), to_signed(16#1ED11#, 20), to_signed(16#1ED6A#, 20),
                                                                              to_signed(16#1EDC2#, 20), to_signed(16#1EE1A#, 20), to_signed(16#1EE72#, 20), to_signed(16#1EECA#, 20),
                                                                              to_signed(16#1EF22#, 20), to_signed(16#1EF7A#, 20), to_signed(16#1EFD2#, 20), to_signed(16#1F02A#, 20),
                                                                              to_signed(16#1F082#, 20), to_signed(16#1F0D9#, 20), to_signed(16#1F131#, 20), to_signed(16#1F189#, 20),
                                                                              to_signed(16#1F1E1#, 20), to_signed(16#1F239#, 20), to_signed(16#1F291#, 20), to_signed(16#1F2E9#, 20),
                                                                              to_signed(16#1F340#, 20), to_signed(16#1F398#, 20), to_signed(16#1F3F0#, 20), to_signed(16#1F448#, 20),
                                                                              to_signed(16#1F49F#, 20), to_signed(16#1F4F7#, 20), to_signed(16#1F54F#, 20), to_signed(16#1F5A6#, 20),
                                                                              to_signed(16#1F5FE#, 20), to_signed(16#1F656#, 20), to_signed(16#1F6AD#, 20), to_signed(16#1F705#, 20),
                                                                              to_signed(16#1F75C#, 20), to_signed(16#1F7B4#, 20), to_signed(16#1F80B#, 20), to_signed(16#1F863#, 20),
                                                                              to_signed(16#1F8BA#, 20), to_signed(16#1F912#, 20), to_signed(16#1F969#, 20), to_signed(16#1F9C1#, 20),
                                                                              to_signed(16#1FA18#, 20), to_signed(16#1FA6F#, 20), to_signed(16#1FAC7#, 20), to_signed(16#1FB1E#, 20),
                                                                              to_signed(16#1FB75#, 20), to_signed(16#1FBCD#, 20), to_signed(16#1FC24#, 20), to_signed(16#1FC7B#, 20),
                                                                              to_signed(16#1FCD3#, 20), to_signed(16#1FD2A#, 20), to_signed(16#1FD81#, 20), to_signed(16#1FDD8#, 20),
                                                                              to_signed(16#1FE2F#, 20), to_signed(16#1FE87#, 20), to_signed(16#1FEDE#, 20), to_signed(16#1FF35#, 20),
                                                                              to_signed(16#1FF8C#, 20), to_signed(16#1FFE3#, 20), to_signed(16#2003A#, 20), to_signed(16#20091#, 20),
                                                                              to_signed(16#200E8#, 20), to_signed(16#2013F#, 20), to_signed(16#20196#, 20), to_signed(16#201ED#, 20),
                                                                              to_signed(16#20244#, 20), to_signed(16#2029B#, 20), to_signed(16#202F2#, 20), to_signed(16#20349#, 20),
                                                                              to_signed(16#203A0#, 20), to_signed(16#203F6#, 20), to_signed(16#2044D#, 20), to_signed(16#204A4#, 20),
                                                                              to_signed(16#204FB#, 20), to_signed(16#20552#, 20), to_signed(16#205A8#, 20), to_signed(16#205FF#, 20),
                                                                              to_signed(16#20656#, 20), to_signed(16#206AC#, 20), to_signed(16#20703#, 20), to_signed(16#2075A#, 20),
                                                                              to_signed(16#207B0#, 20), to_signed(16#20807#, 20), to_signed(16#2085E#, 20), to_signed(16#208B4#, 20),
                                                                              to_signed(16#2090B#, 20), to_signed(16#20961#, 20), to_signed(16#209B8#, 20), to_signed(16#20A0E#, 20),
                                                                              to_signed(16#20A65#, 20), to_signed(16#20ABB#, 20), to_signed(16#20B12#, 20), to_signed(16#20B68#, 20),
                                                                              to_signed(16#20BBE#, 20), to_signed(16#20C15#, 20), to_signed(16#20C6B#, 20), to_signed(16#20CC2#, 20),
                                                                              to_signed(16#20D18#, 20), to_signed(16#20D6E#, 20), to_signed(16#20DC4#, 20), to_signed(16#20E1B#, 20),
                                                                              to_signed(16#20E71#, 20), to_signed(16#20EC7#, 20), to_signed(16#20F1D#, 20), to_signed(16#20F74#, 20),
                                                                              to_signed(16#20FCA#, 20), to_signed(16#21020#, 20), to_signed(16#21076#, 20), to_signed(16#210CC#, 20),
                                                                              to_signed(16#21122#, 20), to_signed(16#21178#, 20), to_signed(16#211CE#, 20), to_signed(16#21224#, 20),
                                                                              to_signed(16#2127A#, 20), to_signed(16#212D0#, 20), to_signed(16#21326#, 20), to_signed(16#2137C#, 20),
                                                                              to_signed(16#213D2#, 20), to_signed(16#21428#, 20), to_signed(16#2147E#, 20), to_signed(16#214D4#, 20),
                                                                              to_signed(16#2152A#, 20), to_signed(16#2157F#, 20), to_signed(16#215D5#, 20), to_signed(16#2162B#, 20),
                                                                              to_signed(16#21681#, 20), to_signed(16#216D6#, 20), to_signed(16#2172C#, 20), to_signed(16#21782#, 20),
                                                                              to_signed(16#217D8#, 20), to_signed(16#2182D#, 20), to_signed(16#21883#, 20), to_signed(16#218D8#, 20),
                                                                              to_signed(16#2192E#, 20), to_signed(16#21984#, 20), to_signed(16#219D9#, 20), to_signed(16#21A2F#, 20),
                                                                              to_signed(16#21A84#, 20), to_signed(16#21ADA#, 20), to_signed(16#21B2F#, 20), to_signed(16#21B85#, 20),
                                                                              to_signed(16#21BDA#, 20), to_signed(16#21C30#, 20), to_signed(16#21C85#, 20), to_signed(16#21CDA#, 20),
                                                                              to_signed(16#21D30#, 20), to_signed(16#21D85#, 20), to_signed(16#21DDA#, 20), to_signed(16#21E30#, 20),
                                                                              to_signed(16#21E85#, 20), to_signed(16#21EDA#, 20), to_signed(16#21F2F#, 20), to_signed(16#21F85#, 20),
                                                                              to_signed(16#21FDA#, 20), to_signed(16#2202F#, 20), to_signed(16#22084#, 20), to_signed(16#220D9#, 20),
                                                                              to_signed(16#2212E#, 20), to_signed(16#22183#, 20), to_signed(16#221D8#, 20), to_signed(16#2222D#, 20),
                                                                              to_signed(16#22283#, 20), to_signed(16#222D8#, 20), to_signed(16#2232D#, 20), to_signed(16#22381#, 20),
                                                                              to_signed(16#223D6#, 20), to_signed(16#2242B#, 20), to_signed(16#22480#, 20), to_signed(16#224D5#, 20),
                                                                              to_signed(16#2252A#, 20), to_signed(16#2257F#, 20), to_signed(16#225D4#, 20), to_signed(16#22628#, 20),
                                                                              to_signed(16#2267D#, 20), to_signed(16#226D2#, 20), to_signed(16#22727#, 20), to_signed(16#2277B#, 20),
                                                                              to_signed(16#227D0#, 20), to_signed(16#22825#, 20), to_signed(16#22879#, 20), to_signed(16#228CE#, 20),
                                                                              to_signed(16#22923#, 20), to_signed(16#22977#, 20), to_signed(16#229CC#, 20), to_signed(16#22A20#, 20),
                                                                              to_signed(16#22A75#, 20), to_signed(16#22AC9#, 20), to_signed(16#22B1E#, 20), to_signed(16#22B72#, 20),
                                                                              to_signed(16#22BC7#, 20), to_signed(16#22C1B#, 20), to_signed(16#22C70#, 20), to_signed(16#22CC4#, 20),
                                                                              to_signed(16#22D18#, 20), to_signed(16#22D6D#, 20), to_signed(16#22DC1#, 20), to_signed(16#22E15#, 20),
                                                                              to_signed(16#22E6A#, 20), to_signed(16#22EBE#, 20), to_signed(16#22F12#, 20), to_signed(16#22F66#, 20),
                                                                              to_signed(16#22FBB#, 20), to_signed(16#2300F#, 20), to_signed(16#23063#, 20), to_signed(16#230B7#, 20),
                                                                              to_signed(16#2310B#, 20), to_signed(16#2315F#, 20), to_signed(16#231B3#, 20), to_signed(16#23207#, 20),
                                                                              to_signed(16#2325B#, 20), to_signed(16#232AF#, 20), to_signed(16#23303#, 20), to_signed(16#23357#, 20),
                                                                              to_signed(16#233AB#, 20), to_signed(16#233FF#, 20), to_signed(16#23453#, 20), to_signed(16#234A7#, 20),
                                                                              to_signed(16#234FB#, 20), to_signed(16#2354F#, 20), to_signed(16#235A2#, 20), to_signed(16#235F6#, 20),
                                                                              to_signed(16#2364A#, 20), to_signed(16#2369E#, 20), to_signed(16#236F1#, 20), to_signed(16#23745#, 20),
                                                                              to_signed(16#23799#, 20), to_signed(16#237ED#, 20), to_signed(16#23840#, 20), to_signed(16#23894#, 20),
                                                                              to_signed(16#238E7#, 20), to_signed(16#2393B#, 20), to_signed(16#2398F#, 20), to_signed(16#239E2#, 20),
                                                                              to_signed(16#23A36#, 20), to_signed(16#23A89#, 20), to_signed(16#23ADD#, 20), to_signed(16#23B30#, 20),
                                                                              to_signed(16#23B83#, 20), to_signed(16#23BD7#, 20), to_signed(16#23C2A#, 20), to_signed(16#23C7E#, 20),
                                                                              to_signed(16#23CD1#, 20), to_signed(16#23D24#, 20), to_signed(16#23D78#, 20), to_signed(16#23DCB#, 20),
                                                                              to_signed(16#23E1E#, 20), to_signed(16#23E71#, 20), to_signed(16#23EC5#, 20), to_signed(16#23F18#, 20),
                                                                              to_signed(16#23F6B#, 20), to_signed(16#23FBE#, 20), to_signed(16#24011#, 20), to_signed(16#24064#, 20),
                                                                              to_signed(16#240B7#, 20), to_signed(16#2410A#, 20), to_signed(16#2415D#, 20), to_signed(16#241B0#, 20),
                                                                              to_signed(16#24203#, 20), to_signed(16#24256#, 20), to_signed(16#242A9#, 20), to_signed(16#242FC#, 20),
                                                                              to_signed(16#2434F#, 20), to_signed(16#243A2#, 20), to_signed(16#243F5#, 20), to_signed(16#24448#, 20),
                                                                              to_signed(16#2449B#, 20), to_signed(16#244ED#, 20), to_signed(16#24540#, 20), to_signed(16#24593#, 20),
                                                                              to_signed(16#245E6#, 20), to_signed(16#24638#, 20), to_signed(16#2468B#, 20), to_signed(16#246DE#, 20),
                                                                              to_signed(16#24730#, 20), to_signed(16#24783#, 20), to_signed(16#247D6#, 20), to_signed(16#24828#, 20),
                                                                              to_signed(16#2487B#, 20), to_signed(16#248CD#, 20), to_signed(16#24920#, 20), to_signed(16#24972#, 20),
                                                                              to_signed(16#249C5#, 20), to_signed(16#24A17#, 20), to_signed(16#24A6A#, 20), to_signed(16#24ABC#, 20),
                                                                              to_signed(16#24B0E#, 20), to_signed(16#24B61#, 20), to_signed(16#24BB3#, 20), to_signed(16#24C05#, 20),
                                                                              to_signed(16#24C58#, 20), to_signed(16#24CAA#, 20), to_signed(16#24CFC#, 20), to_signed(16#24D4E#, 20),
                                                                              to_signed(16#24DA1#, 20), to_signed(16#24DF3#, 20), to_signed(16#24E45#, 20), to_signed(16#24E97#, 20),
                                                                              to_signed(16#24EE9#, 20), to_signed(16#24F3B#, 20), to_signed(16#24F8D#, 20), to_signed(16#24FDF#, 20),
                                                                              to_signed(16#25031#, 20), to_signed(16#25083#, 20), to_signed(16#250D5#, 20), to_signed(16#25127#, 20),
                                                                              to_signed(16#25179#, 20), to_signed(16#251CB#, 20), to_signed(16#2521D#, 20), to_signed(16#2526F#, 20),
                                                                              to_signed(16#252C1#, 20), to_signed(16#25313#, 20), to_signed(16#25365#, 20), to_signed(16#253B6#, 20),
                                                                              to_signed(16#25408#, 20), to_signed(16#2545A#, 20), to_signed(16#254AC#, 20), to_signed(16#254FD#, 20),
                                                                              to_signed(16#2554F#, 20), to_signed(16#255A1#, 20), to_signed(16#255F2#, 20), to_signed(16#25644#, 20),
                                                                              to_signed(16#25695#, 20), to_signed(16#256E7#, 20), to_signed(16#25738#, 20), to_signed(16#2578A#, 20),
                                                                              to_signed(16#257DB#, 20), to_signed(16#2582D#, 20), to_signed(16#2587E#, 20), to_signed(16#258D0#, 20),
                                                                              to_signed(16#25921#, 20), to_signed(16#25972#, 20), to_signed(16#259C4#, 20), to_signed(16#25A15#, 20),
                                                                              to_signed(16#25A66#, 20), to_signed(16#25AB8#, 20), to_signed(16#25B09#, 20), to_signed(16#25B5A#, 20),
                                                                              to_signed(16#25BAB#, 20), to_signed(16#25BFD#, 20), to_signed(16#25C4E#, 20), to_signed(16#25C9F#, 20),
                                                                              to_signed(16#25CF0#, 20), to_signed(16#25D41#, 20), to_signed(16#25D92#, 20), to_signed(16#25DE3#, 20),
                                                                              to_signed(16#25E34#, 20), to_signed(16#25E85#, 20), to_signed(16#25ED6#, 20), to_signed(16#25F27#, 20),
                                                                              to_signed(16#25F78#, 20), to_signed(16#25FC9#, 20), to_signed(16#2601A#, 20), to_signed(16#2606B#, 20),
                                                                              to_signed(16#260BC#, 20), to_signed(16#2610D#, 20), to_signed(16#2615D#, 20), to_signed(16#261AE#, 20),
                                                                              to_signed(16#261FF#, 20), to_signed(16#26250#, 20), to_signed(16#262A0#, 20), to_signed(16#262F1#, 20),
                                                                              to_signed(16#26342#, 20), to_signed(16#26392#, 20), to_signed(16#263E3#, 20), to_signed(16#26434#, 20),
                                                                              to_signed(16#26484#, 20), to_signed(16#264D5#, 20), to_signed(16#26525#, 20), to_signed(16#26576#, 20),
                                                                              to_signed(16#265C6#, 20), to_signed(16#26617#, 20), to_signed(16#26667#, 20), to_signed(16#266B8#, 20),
                                                                              to_signed(16#26708#, 20), to_signed(16#26758#, 20), to_signed(16#267A9#, 20), to_signed(16#267F9#, 20),
                                                                              to_signed(16#26849#, 20), to_signed(16#2689A#, 20), to_signed(16#268EA#, 20), to_signed(16#2693A#, 20),
                                                                              to_signed(16#2698A#, 20), to_signed(16#269DA#, 20), to_signed(16#26A2B#, 20), to_signed(16#26A7B#, 20),
                                                                              to_signed(16#26ACB#, 20), to_signed(16#26B1B#, 20), to_signed(16#26B6B#, 20), to_signed(16#26BBB#, 20),
                                                                              to_signed(16#26C0B#, 20), to_signed(16#26C5B#, 20), to_signed(16#26CAB#, 20), to_signed(16#26CFB#, 20),
                                                                              to_signed(16#26D4B#, 20), to_signed(16#26D9B#, 20), to_signed(16#26DEB#, 20), to_signed(16#26E3B#, 20),
                                                                              to_signed(16#26E8A#, 20), to_signed(16#26EDA#, 20), to_signed(16#26F2A#, 20), to_signed(16#26F7A#, 20),
                                                                              to_signed(16#26FC9#, 20), to_signed(16#27019#, 20), to_signed(16#27069#, 20), to_signed(16#270B9#, 20),
                                                                              to_signed(16#27108#, 20), to_signed(16#27158#, 20), to_signed(16#271A7#, 20), to_signed(16#271F7#, 20),
                                                                              to_signed(16#27247#, 20), to_signed(16#27296#, 20), to_signed(16#272E6#, 20), to_signed(16#27335#, 20),
                                                                              to_signed(16#27384#, 20), to_signed(16#273D4#, 20), to_signed(16#27423#, 20), to_signed(16#27473#, 20),
                                                                              to_signed(16#274C2#, 20), to_signed(16#27511#, 20), to_signed(16#27561#, 20), to_signed(16#275B0#, 20),
                                                                              to_signed(16#275FF#, 20), to_signed(16#2764F#, 20), to_signed(16#2769E#, 20), to_signed(16#276ED#, 20),
                                                                              to_signed(16#2773C#, 20), to_signed(16#2778B#, 20), to_signed(16#277DA#, 20), to_signed(16#27829#, 20),
                                                                              to_signed(16#27879#, 20), to_signed(16#278C8#, 20), to_signed(16#27917#, 20), to_signed(16#27966#, 20),
                                                                              to_signed(16#279B5#, 20), to_signed(16#27A04#, 20), to_signed(16#27A52#, 20), to_signed(16#27AA1#, 20),
                                                                              to_signed(16#27AF0#, 20), to_signed(16#27B3F#, 20), to_signed(16#27B8E#, 20), to_signed(16#27BDD#, 20),
                                                                              to_signed(16#27C2C#, 20), to_signed(16#27C7A#, 20), to_signed(16#27CC9#, 20), to_signed(16#27D18#, 20),
                                                                              to_signed(16#27D66#, 20), to_signed(16#27DB5#, 20), to_signed(16#27E04#, 20), to_signed(16#27E52#, 20),
                                                                              to_signed(16#27EA1#, 20), to_signed(16#27EF0#, 20), to_signed(16#27F3E#, 20), to_signed(16#27F8D#, 20),
                                                                              to_signed(16#27FDB#, 20), to_signed(16#2802A#, 20), to_signed(16#28078#, 20), to_signed(16#280C7#, 20),
                                                                              to_signed(16#28115#, 20), to_signed(16#28163#, 20), to_signed(16#281B2#, 20), to_signed(16#28200#, 20),
                                                                              to_signed(16#2824E#, 20), to_signed(16#2829D#, 20), to_signed(16#282EB#, 20), to_signed(16#28339#, 20),
                                                                              to_signed(16#28387#, 20), to_signed(16#283D5#, 20), to_signed(16#28424#, 20), to_signed(16#28472#, 20),
                                                                              to_signed(16#284C0#, 20), to_signed(16#2850E#, 20), to_signed(16#2855C#, 20), to_signed(16#285AA#, 20),
                                                                              to_signed(16#285F8#, 20), to_signed(16#28646#, 20), to_signed(16#28694#, 20), to_signed(16#286E2#, 20),
                                                                              to_signed(16#28730#, 20), to_signed(16#2877E#, 20), to_signed(16#287CC#, 20), to_signed(16#2881A#, 20),
                                                                              to_signed(16#28867#, 20), to_signed(16#288B5#, 20), to_signed(16#28903#, 20), to_signed(16#28951#, 20),
                                                                              to_signed(16#2899E#, 20), to_signed(16#289EC#, 20), to_signed(16#28A3A#, 20), to_signed(16#28A87#, 20),
                                                                              to_signed(16#28AD5#, 20), to_signed(16#28B23#, 20), to_signed(16#28B70#, 20), to_signed(16#28BBE#, 20),
                                                                              to_signed(16#28C0B#, 20), to_signed(16#28C59#, 20), to_signed(16#28CA6#, 20), to_signed(16#28CF4#, 20),
                                                                              to_signed(16#28D41#, 20), to_signed(16#28D8F#, 20), to_signed(16#28DDC#, 20), to_signed(16#28E29#, 20),
                                                                              to_signed(16#28E77#, 20), to_signed(16#28EC4#, 20), to_signed(16#28F11#, 20), to_signed(16#28F5E#, 20),
                                                                              to_signed(16#28FAC#, 20), to_signed(16#28FF9#, 20), to_signed(16#29046#, 20), to_signed(16#29093#, 20),
                                                                              to_signed(16#290E0#, 20), to_signed(16#2912E#, 20), to_signed(16#2917B#, 20), to_signed(16#291C8#, 20),
                                                                              to_signed(16#29215#, 20), to_signed(16#29262#, 20), to_signed(16#292AF#, 20), to_signed(16#292FC#, 20),
                                                                              to_signed(16#29349#, 20), to_signed(16#29395#, 20), to_signed(16#293E2#, 20), to_signed(16#2942F#, 20),
                                                                              to_signed(16#2947C#, 20), to_signed(16#294C9#, 20), to_signed(16#29516#, 20), to_signed(16#29562#, 20),
                                                                              to_signed(16#295AF#, 20), to_signed(16#295FC#, 20), to_signed(16#29649#, 20), to_signed(16#29695#, 20),
                                                                              to_signed(16#296E2#, 20), to_signed(16#2972E#, 20), to_signed(16#2977B#, 20), to_signed(16#297C8#, 20),
                                                                              to_signed(16#29814#, 20), to_signed(16#29861#, 20), to_signed(16#298AD#, 20), to_signed(16#298FA#, 20),
                                                                              to_signed(16#29946#, 20), to_signed(16#29992#, 20), to_signed(16#299DF#, 20), to_signed(16#29A2B#, 20),
                                                                              to_signed(16#29A78#, 20), to_signed(16#29AC4#, 20), to_signed(16#29B10#, 20), to_signed(16#29B5C#, 20),
                                                                              to_signed(16#29BA9#, 20), to_signed(16#29BF5#, 20), to_signed(16#29C41#, 20), to_signed(16#29C8D#, 20),
                                                                              to_signed(16#29CD9#, 20), to_signed(16#29D25#, 20), to_signed(16#29D72#, 20), to_signed(16#29DBE#, 20),
                                                                              to_signed(16#29E0A#, 20), to_signed(16#29E56#, 20), to_signed(16#29EA2#, 20), to_signed(16#29EEE#, 20),
                                                                              to_signed(16#29F3A#, 20), to_signed(16#29F85#, 20), to_signed(16#29FD1#, 20), to_signed(16#2A01D#, 20),
                                                                              to_signed(16#2A069#, 20), to_signed(16#2A0B5#, 20), to_signed(16#2A101#, 20), to_signed(16#2A14C#, 20),
                                                                              to_signed(16#2A198#, 20), to_signed(16#2A1E4#, 20), to_signed(16#2A22F#, 20), to_signed(16#2A27B#, 20),
                                                                              to_signed(16#2A2C7#, 20), to_signed(16#2A312#, 20), to_signed(16#2A35E#, 20), to_signed(16#2A3A9#, 20),
                                                                              to_signed(16#2A3F5#, 20), to_signed(16#2A441#, 20), to_signed(16#2A48C#, 20), to_signed(16#2A4D7#, 20),
                                                                              to_signed(16#2A523#, 20), to_signed(16#2A56E#, 20), to_signed(16#2A5BA#, 20), to_signed(16#2A605#, 20),
                                                                              to_signed(16#2A650#, 20), to_signed(16#2A69C#, 20), to_signed(16#2A6E7#, 20), to_signed(16#2A732#, 20),
                                                                              to_signed(16#2A77D#, 20), to_signed(16#2A7C9#, 20), to_signed(16#2A814#, 20), to_signed(16#2A85F#, 20),
                                                                              to_signed(16#2A8AA#, 20), to_signed(16#2A8F5#, 20), to_signed(16#2A940#, 20), to_signed(16#2A98B#, 20),
                                                                              to_signed(16#2A9D6#, 20), to_signed(16#2AA21#, 20), to_signed(16#2AA6C#, 20), to_signed(16#2AAB7#, 20),
                                                                              to_signed(16#2AB02#, 20), to_signed(16#2AB4D#, 20), to_signed(16#2AB98#, 20), to_signed(16#2ABE3#, 20),
                                                                              to_signed(16#2AC2D#, 20), to_signed(16#2AC78#, 20), to_signed(16#2ACC3#, 20), to_signed(16#2AD0E#, 20),
                                                                              to_signed(16#2AD58#, 20), to_signed(16#2ADA3#, 20), to_signed(16#2ADEE#, 20), to_signed(16#2AE38#, 20),
                                                                              to_signed(16#2AE83#, 20), to_signed(16#2AECE#, 20), to_signed(16#2AF18#, 20), to_signed(16#2AF63#, 20),
                                                                              to_signed(16#2AFAD#, 20), to_signed(16#2AFF8#, 20), to_signed(16#2B042#, 20), to_signed(16#2B08C#, 20),
                                                                              to_signed(16#2B0D7#, 20), to_signed(16#2B121#, 20), to_signed(16#2B16C#, 20), to_signed(16#2B1B6#, 20),
                                                                              to_signed(16#2B200#, 20), to_signed(16#2B24A#, 20), to_signed(16#2B295#, 20), to_signed(16#2B2DF#, 20),
                                                                              to_signed(16#2B329#, 20), to_signed(16#2B373#, 20), to_signed(16#2B3BD#, 20), to_signed(16#2B408#, 20),
                                                                              to_signed(16#2B452#, 20), to_signed(16#2B49C#, 20), to_signed(16#2B4E6#, 20), to_signed(16#2B530#, 20),
                                                                              to_signed(16#2B57A#, 20), to_signed(16#2B5C4#, 20), to_signed(16#2B60E#, 20), to_signed(16#2B658#, 20),
                                                                              to_signed(16#2B6A1#, 20), to_signed(16#2B6EB#, 20), to_signed(16#2B735#, 20), to_signed(16#2B77F#, 20),
                                                                              to_signed(16#2B7C9#, 20), to_signed(16#2B812#, 20), to_signed(16#2B85C#, 20), to_signed(16#2B8A6#, 20),
                                                                              to_signed(16#2B8EF#, 20), to_signed(16#2B939#, 20), to_signed(16#2B983#, 20), to_signed(16#2B9CC#, 20),
                                                                              to_signed(16#2BA16#, 20), to_signed(16#2BA5F#, 20), to_signed(16#2BAA9#, 20), to_signed(16#2BAF2#, 20),
                                                                              to_signed(16#2BB3C#, 20), to_signed(16#2BB85#, 20), to_signed(16#2BBCF#, 20), to_signed(16#2BC18#, 20),
                                                                              to_signed(16#2BC61#, 20), to_signed(16#2BCAB#, 20), to_signed(16#2BCF4#, 20), to_signed(16#2BD3D#, 20),
                                                                              to_signed(16#2BD87#, 20), to_signed(16#2BDD0#, 20), to_signed(16#2BE19#, 20), to_signed(16#2BE62#, 20),
                                                                              to_signed(16#2BEAB#, 20), to_signed(16#2BEF4#, 20), to_signed(16#2BF3D#, 20), to_signed(16#2BF87#, 20),
                                                                              to_signed(16#2BFD0#, 20), to_signed(16#2C019#, 20), to_signed(16#2C062#, 20), to_signed(16#2C0AB#, 20),
                                                                              to_signed(16#2C0F3#, 20), to_signed(16#2C13C#, 20), to_signed(16#2C185#, 20), to_signed(16#2C1CE#, 20),
                                                                              to_signed(16#2C217#, 20), to_signed(16#2C260#, 20), to_signed(16#2C2A8#, 20), to_signed(16#2C2F1#, 20),
                                                                              to_signed(16#2C33A#, 20), to_signed(16#2C383#, 20), to_signed(16#2C3CB#, 20), to_signed(16#2C414#, 20),
                                                                              to_signed(16#2C45D#, 20), to_signed(16#2C4A5#, 20), to_signed(16#2C4EE#, 20), to_signed(16#2C536#, 20),
                                                                              to_signed(16#2C57F#, 20), to_signed(16#2C5C7#, 20), to_signed(16#2C610#, 20), to_signed(16#2C658#, 20),
                                                                              to_signed(16#2C6A0#, 20), to_signed(16#2C6E9#, 20), to_signed(16#2C731#, 20), to_signed(16#2C779#, 20),
                                                                              to_signed(16#2C7C2#, 20), to_signed(16#2C80A#, 20), to_signed(16#2C852#, 20), to_signed(16#2C89A#, 20),
                                                                              to_signed(16#2C8E3#, 20), to_signed(16#2C92B#, 20), to_signed(16#2C973#, 20), to_signed(16#2C9BB#, 20),
                                                                              to_signed(16#2CA03#, 20), to_signed(16#2CA4B#, 20), to_signed(16#2CA93#, 20), to_signed(16#2CADB#, 20),
                                                                              to_signed(16#2CB23#, 20), to_signed(16#2CB6B#, 20), to_signed(16#2CBB3#, 20), to_signed(16#2CBFB#, 20),
                                                                              to_signed(16#2CC43#, 20), to_signed(16#2CC8B#, 20), to_signed(16#2CCD2#, 20), to_signed(16#2CD1A#, 20),
                                                                              to_signed(16#2CD62#, 20), to_signed(16#2CDAA#, 20), to_signed(16#2CDF1#, 20), to_signed(16#2CE39#, 20),
                                                                              to_signed(16#2CE81#, 20), to_signed(16#2CEC8#, 20), to_signed(16#2CF10#, 20), to_signed(16#2CF57#, 20),
                                                                              to_signed(16#2CF9F#, 20), to_signed(16#2CFE6#, 20), to_signed(16#2D02E#, 20), to_signed(16#2D075#, 20),
                                                                              to_signed(16#2D0BD#, 20), to_signed(16#2D104#, 20), to_signed(16#2D14C#, 20), to_signed(16#2D193#, 20),
                                                                              to_signed(16#2D1DA#, 20), to_signed(16#2D222#, 20), to_signed(16#2D269#, 20), to_signed(16#2D2B0#, 20),
                                                                              to_signed(16#2D2F7#, 20), to_signed(16#2D33E#, 20), to_signed(16#2D386#, 20), to_signed(16#2D3CD#, 20),
                                                                              to_signed(16#2D414#, 20), to_signed(16#2D45B#, 20), to_signed(16#2D4A2#, 20), to_signed(16#2D4E9#, 20),
                                                                              to_signed(16#2D530#, 20), to_signed(16#2D577#, 20), to_signed(16#2D5BE#, 20), to_signed(16#2D605#, 20),
                                                                              to_signed(16#2D64C#, 20), to_signed(16#2D692#, 20), to_signed(16#2D6D9#, 20), to_signed(16#2D720#, 20),
                                                                              to_signed(16#2D767#, 20), to_signed(16#2D7AE#, 20), to_signed(16#2D7F4#, 20), to_signed(16#2D83B#, 20),
                                                                              to_signed(16#2D882#, 20), to_signed(16#2D8C8#, 20), to_signed(16#2D90F#, 20), to_signed(16#2D956#, 20),
                                                                              to_signed(16#2D99C#, 20), to_signed(16#2D9E3#, 20), to_signed(16#2DA29#, 20), to_signed(16#2DA70#, 20),
                                                                              to_signed(16#2DAB6#, 20), to_signed(16#2DAFC#, 20), to_signed(16#2DB43#, 20), to_signed(16#2DB89#, 20),
                                                                              to_signed(16#2DBCF#, 20), to_signed(16#2DC16#, 20), to_signed(16#2DC5C#, 20), to_signed(16#2DCA2#, 20),
                                                                              to_signed(16#2DCE9#, 20), to_signed(16#2DD2F#, 20), to_signed(16#2DD75#, 20), to_signed(16#2DDBB#, 20),
                                                                              to_signed(16#2DE01#, 20), to_signed(16#2DE47#, 20), to_signed(16#2DE8D#, 20), to_signed(16#2DED3#, 20),
                                                                              to_signed(16#2DF19#, 20), to_signed(16#2DF5F#, 20), to_signed(16#2DFA5#, 20), to_signed(16#2DFEB#, 20),
                                                                              to_signed(16#2E031#, 20), to_signed(16#2E077#, 20), to_signed(16#2E0BD#, 20), to_signed(16#2E103#, 20),
                                                                              to_signed(16#2E148#, 20), to_signed(16#2E18E#, 20), to_signed(16#2E1D4#, 20), to_signed(16#2E21A#, 20),
                                                                              to_signed(16#2E25F#, 20), to_signed(16#2E2A5#, 20), to_signed(16#2E2EA#, 20), to_signed(16#2E330#, 20),
                                                                              to_signed(16#2E376#, 20), to_signed(16#2E3BB#, 20), to_signed(16#2E401#, 20), to_signed(16#2E446#, 20),
                                                                              to_signed(16#2E48C#, 20), to_signed(16#2E4D1#, 20), to_signed(16#2E516#, 20), to_signed(16#2E55C#, 20),
                                                                              to_signed(16#2E5A1#, 20), to_signed(16#2E5E6#, 20), to_signed(16#2E62C#, 20), to_signed(16#2E671#, 20),
                                                                              to_signed(16#2E6B6#, 20), to_signed(16#2E6FB#, 20), to_signed(16#2E740#, 20), to_signed(16#2E786#, 20),
                                                                              to_signed(16#2E7CB#, 20), to_signed(16#2E810#, 20), to_signed(16#2E855#, 20), to_signed(16#2E89A#, 20),
                                                                              to_signed(16#2E8DF#, 20), to_signed(16#2E924#, 20), to_signed(16#2E969#, 20), to_signed(16#2E9AE#, 20),
                                                                              to_signed(16#2E9F3#, 20), to_signed(16#2EA37#, 20), to_signed(16#2EA7C#, 20), to_signed(16#2EAC1#, 20),
                                                                              to_signed(16#2EB06#, 20), to_signed(16#2EB4B#, 20), to_signed(16#2EB8F#, 20), to_signed(16#2EBD4#, 20),
                                                                              to_signed(16#2EC19#, 20), to_signed(16#2EC5D#, 20), to_signed(16#2ECA2#, 20), to_signed(16#2ECE6#, 20),
                                                                              to_signed(16#2ED2B#, 20), to_signed(16#2ED70#, 20), to_signed(16#2EDB4#, 20), to_signed(16#2EDF8#, 20),
                                                                              to_signed(16#2EE3D#, 20), to_signed(16#2EE81#, 20), to_signed(16#2EEC6#, 20), to_signed(16#2EF0A#, 20),
                                                                              to_signed(16#2EF4E#, 20), to_signed(16#2EF93#, 20), to_signed(16#2EFD7#, 20), to_signed(16#2F01B#, 20),
                                                                              to_signed(16#2F05F#, 20), to_signed(16#2F0A4#, 20), to_signed(16#2F0E8#, 20), to_signed(16#2F12C#, 20),
                                                                              to_signed(16#2F170#, 20), to_signed(16#2F1B4#, 20), to_signed(16#2F1F8#, 20), to_signed(16#2F23C#, 20),
                                                                              to_signed(16#2F280#, 20), to_signed(16#2F2C4#, 20), to_signed(16#2F308#, 20), to_signed(16#2F34C#, 20),
                                                                              to_signed(16#2F390#, 20), to_signed(16#2F3D4#, 20), to_signed(16#2F417#, 20), to_signed(16#2F45B#, 20),
                                                                              to_signed(16#2F49F#, 20), to_signed(16#2F4E3#, 20), to_signed(16#2F526#, 20), to_signed(16#2F56A#, 20),
                                                                              to_signed(16#2F5AE#, 20), to_signed(16#2F5F1#, 20), to_signed(16#2F635#, 20), to_signed(16#2F678#, 20),
                                                                              to_signed(16#2F6BC#, 20), to_signed(16#2F6FF#, 20), to_signed(16#2F743#, 20), to_signed(16#2F786#, 20),
                                                                              to_signed(16#2F7CA#, 20), to_signed(16#2F80D#, 20), to_signed(16#2F850#, 20), to_signed(16#2F894#, 20),
                                                                              to_signed(16#2F8D7#, 20), to_signed(16#2F91A#, 20), to_signed(16#2F95E#, 20), to_signed(16#2F9A1#, 20),
                                                                              to_signed(16#2F9E4#, 20), to_signed(16#2FA27#, 20), to_signed(16#2FA6A#, 20), to_signed(16#2FAAD#, 20),
                                                                              to_signed(16#2FAF0#, 20), to_signed(16#2FB33#, 20), to_signed(16#2FB76#, 20), to_signed(16#2FBB9#, 20),
                                                                              to_signed(16#2FBFC#, 20), to_signed(16#2FC3F#, 20), to_signed(16#2FC82#, 20), to_signed(16#2FCC5#, 20),
                                                                              to_signed(16#2FD08#, 20), to_signed(16#2FD4B#, 20), to_signed(16#2FD8E#, 20), to_signed(16#2FDD0#, 20),
                                                                              to_signed(16#2FE13#, 20), to_signed(16#2FE56#, 20), to_signed(16#2FE98#, 20), to_signed(16#2FEDB#, 20),
                                                                              to_signed(16#2FF1E#, 20), to_signed(16#2FF60#, 20), to_signed(16#2FFA3#, 20), to_signed(16#2FFE5#, 20),
                                                                              to_signed(16#30028#, 20), to_signed(16#3006A#, 20), to_signed(16#300AD#, 20), to_signed(16#300EF#, 20),
                                                                              to_signed(16#30131#, 20), to_signed(16#30174#, 20), to_signed(16#301B6#, 20), to_signed(16#301F8#, 20),
                                                                              to_signed(16#3023B#, 20), to_signed(16#3027D#, 20), to_signed(16#302BF#, 20), to_signed(16#30301#, 20),
                                                                              to_signed(16#30343#, 20), to_signed(16#30386#, 20), to_signed(16#303C8#, 20), to_signed(16#3040A#, 20),
                                                                              to_signed(16#3044C#, 20), to_signed(16#3048E#, 20), to_signed(16#304D0#, 20), to_signed(16#30512#, 20),
                                                                              to_signed(16#30554#, 20), to_signed(16#30595#, 20), to_signed(16#305D7#, 20), to_signed(16#30619#, 20),
                                                                              to_signed(16#3065B#, 20), to_signed(16#3069D#, 20), to_signed(16#306DE#, 20), to_signed(16#30720#, 20),
                                                                              to_signed(16#30762#, 20), to_signed(16#307A3#, 20), to_signed(16#307E5#, 20), to_signed(16#30827#, 20),
                                                                              to_signed(16#30868#, 20), to_signed(16#308AA#, 20), to_signed(16#308EB#, 20), to_signed(16#3092D#, 20),
                                                                              to_signed(16#3096E#, 20), to_signed(16#309B0#, 20), to_signed(16#309F1#, 20), to_signed(16#30A32#, 20),
                                                                              to_signed(16#30A74#, 20), to_signed(16#30AB5#, 20), to_signed(16#30AF6#, 20), to_signed(16#30B37#, 20),
                                                                              to_signed(16#30B79#, 20), to_signed(16#30BBA#, 20), to_signed(16#30BFB#, 20), to_signed(16#30C3C#, 20),
                                                                              to_signed(16#30C7D#, 20), to_signed(16#30CBE#, 20), to_signed(16#30CFF#, 20), to_signed(16#30D40#, 20),
                                                                              to_signed(16#30D81#, 20), to_signed(16#30DC2#, 20), to_signed(16#30E03#, 20), to_signed(16#30E44#, 20),
                                                                              to_signed(16#30E85#, 20), to_signed(16#30EC6#, 20), to_signed(16#30F06#, 20), to_signed(16#30F47#, 20),
                                                                              to_signed(16#30F88#, 20), to_signed(16#30FC9#, 20), to_signed(16#31009#, 20), to_signed(16#3104A#, 20),
                                                                              to_signed(16#3108B#, 20), to_signed(16#310CB#, 20), to_signed(16#3110C#, 20), to_signed(16#3114C#, 20),
                                                                              to_signed(16#3118D#, 20), to_signed(16#311CD#, 20), to_signed(16#3120E#, 20), to_signed(16#3124E#, 20),
                                                                              to_signed(16#3128F#, 20), to_signed(16#312CF#, 20), to_signed(16#3130F#, 20), to_signed(16#31350#, 20),
                                                                              to_signed(16#31390#, 20), to_signed(16#313D0#, 20), to_signed(16#31410#, 20), to_signed(16#31450#, 20),
                                                                              to_signed(16#31491#, 20), to_signed(16#314D1#, 20), to_signed(16#31511#, 20), to_signed(16#31551#, 20),
                                                                              to_signed(16#31591#, 20), to_signed(16#315D1#, 20), to_signed(16#31611#, 20), to_signed(16#31651#, 20),
                                                                              to_signed(16#31691#, 20), to_signed(16#316D1#, 20), to_signed(16#31710#, 20), to_signed(16#31750#, 20),
                                                                              to_signed(16#31790#, 20), to_signed(16#317D0#, 20), to_signed(16#31810#, 20), to_signed(16#3184F#, 20),
                                                                              to_signed(16#3188F#, 20), to_signed(16#318CF#, 20), to_signed(16#3190E#, 20), to_signed(16#3194E#, 20),
                                                                              to_signed(16#3198D#, 20), to_signed(16#319CD#, 20), to_signed(16#31A0C#, 20), to_signed(16#31A4C#, 20),
                                                                              to_signed(16#31A8B#, 20), to_signed(16#31ACB#, 20), to_signed(16#31B0A#, 20), to_signed(16#31B49#, 20),
                                                                              to_signed(16#31B89#, 20), to_signed(16#31BC8#, 20), to_signed(16#31C07#, 20), to_signed(16#31C46#, 20),
                                                                              to_signed(16#31C86#, 20), to_signed(16#31CC5#, 20), to_signed(16#31D04#, 20), to_signed(16#31D43#, 20),
                                                                              to_signed(16#31D82#, 20), to_signed(16#31DC1#, 20), to_signed(16#31E00#, 20), to_signed(16#31E3F#, 20),
                                                                              to_signed(16#31E7E#, 20), to_signed(16#31EBD#, 20), to_signed(16#31EFC#, 20), to_signed(16#31F3B#, 20),
                                                                              to_signed(16#31F7A#, 20), to_signed(16#31FB8#, 20), to_signed(16#31FF7#, 20), to_signed(16#32036#, 20),
                                                                              to_signed(16#32075#, 20), to_signed(16#320B3#, 20), to_signed(16#320F2#, 20), to_signed(16#32131#, 20),
                                                                              to_signed(16#3216F#, 20), to_signed(16#321AE#, 20), to_signed(16#321EC#, 20), to_signed(16#3222B#, 20),
                                                                              to_signed(16#32269#, 20), to_signed(16#322A8#, 20), to_signed(16#322E6#, 20), to_signed(16#32324#, 20),
                                                                              to_signed(16#32363#, 20), to_signed(16#323A1#, 20), to_signed(16#323DF#, 20), to_signed(16#3241E#, 20),
                                                                              to_signed(16#3245C#, 20), to_signed(16#3249A#, 20), to_signed(16#324D8#, 20), to_signed(16#32516#, 20),
                                                                              to_signed(16#32555#, 20), to_signed(16#32593#, 20), to_signed(16#325D1#, 20), to_signed(16#3260F#, 20),
                                                                              to_signed(16#3264D#, 20), to_signed(16#3268B#, 20), to_signed(16#326C9#, 20), to_signed(16#32706#, 20),
                                                                              to_signed(16#32744#, 20), to_signed(16#32782#, 20), to_signed(16#327C0#, 20), to_signed(16#327FE#, 20),
                                                                              to_signed(16#3283B#, 20), to_signed(16#32879#, 20), to_signed(16#328B7#, 20), to_signed(16#328F4#, 20),
                                                                              to_signed(16#32932#, 20), to_signed(16#32970#, 20), to_signed(16#329AD#, 20), to_signed(16#329EB#, 20),
                                                                              to_signed(16#32A28#, 20), to_signed(16#32A66#, 20), to_signed(16#32AA3#, 20), to_signed(16#32AE1#, 20),
                                                                              to_signed(16#32B1E#, 20), to_signed(16#32B5B#, 20), to_signed(16#32B99#, 20), to_signed(16#32BD6#, 20),
                                                                              to_signed(16#32C13#, 20), to_signed(16#32C50#, 20), to_signed(16#32C8E#, 20), to_signed(16#32CCB#, 20),
                                                                              to_signed(16#32D08#, 20), to_signed(16#32D45#, 20), to_signed(16#32D82#, 20), to_signed(16#32DBF#, 20),
                                                                              to_signed(16#32DFC#, 20), to_signed(16#32E39#, 20), to_signed(16#32E76#, 20), to_signed(16#32EB3#, 20),
                                                                              to_signed(16#32EF0#, 20), to_signed(16#32F2D#, 20), to_signed(16#32F6A#, 20), to_signed(16#32FA6#, 20),
                                                                              to_signed(16#32FE3#, 20), to_signed(16#33020#, 20), to_signed(16#3305D#, 20), to_signed(16#33099#, 20),
                                                                              to_signed(16#330D6#, 20), to_signed(16#33112#, 20), to_signed(16#3314F#, 20), to_signed(16#3318C#, 20),
                                                                              to_signed(16#331C8#, 20), to_signed(16#33205#, 20), to_signed(16#33241#, 20), to_signed(16#3327E#, 20),
                                                                              to_signed(16#332BA#, 20), to_signed(16#332F6#, 20), to_signed(16#33333#, 20), to_signed(16#3336F#, 20),
                                                                              to_signed(16#333AB#, 20), to_signed(16#333E7#, 20), to_signed(16#33424#, 20), to_signed(16#33460#, 20),
                                                                              to_signed(16#3349C#, 20), to_signed(16#334D8#, 20), to_signed(16#33514#, 20), to_signed(16#33550#, 20),
                                                                              to_signed(16#3358C#, 20), to_signed(16#335C8#, 20), to_signed(16#33604#, 20), to_signed(16#33640#, 20),
                                                                              to_signed(16#3367C#, 20), to_signed(16#336B8#, 20), to_signed(16#336F4#, 20), to_signed(16#33730#, 20),
                                                                              to_signed(16#3376B#, 20), to_signed(16#337A7#, 20), to_signed(16#337E3#, 20), to_signed(16#3381E#, 20),
                                                                              to_signed(16#3385A#, 20), to_signed(16#33896#, 20), to_signed(16#338D1#, 20), to_signed(16#3390D#, 20),
                                                                              to_signed(16#33948#, 20), to_signed(16#33984#, 20), to_signed(16#339BF#, 20), to_signed(16#339FB#, 20),
                                                                              to_signed(16#33A36#, 20), to_signed(16#33A72#, 20), to_signed(16#33AAD#, 20), to_signed(16#33AE8#, 20),
                                                                              to_signed(16#33B24#, 20), to_signed(16#33B5F#, 20), to_signed(16#33B9A#, 20), to_signed(16#33BD5#, 20),
                                                                              to_signed(16#33C10#, 20), to_signed(16#33C4B#, 20), to_signed(16#33C87#, 20), to_signed(16#33CC2#, 20),
                                                                              to_signed(16#33CFD#, 20), to_signed(16#33D38#, 20), to_signed(16#33D73#, 20), to_signed(16#33DAE#, 20),
                                                                              to_signed(16#33DE8#, 20), to_signed(16#33E23#, 20), to_signed(16#33E5E#, 20), to_signed(16#33E99#, 20),
                                                                              to_signed(16#33ED4#, 20), to_signed(16#33F0F#, 20), to_signed(16#33F49#, 20), to_signed(16#33F84#, 20),
                                                                              to_signed(16#33FBF#, 20), to_signed(16#33FF9#, 20), to_signed(16#34034#, 20), to_signed(16#3406E#, 20),
                                                                              to_signed(16#340A9#, 20), to_signed(16#340E3#, 20), to_signed(16#3411E#, 20), to_signed(16#34158#, 20),
                                                                              to_signed(16#34193#, 20), to_signed(16#341CD#, 20), to_signed(16#34207#, 20), to_signed(16#34242#, 20),
                                                                              to_signed(16#3427C#, 20), to_signed(16#342B6#, 20), to_signed(16#342F1#, 20), to_signed(16#3432B#, 20),
                                                                              to_signed(16#34365#, 20), to_signed(16#3439F#, 20), to_signed(16#343D9#, 20), to_signed(16#34413#, 20),
                                                                              to_signed(16#3444D#, 20), to_signed(16#34487#, 20), to_signed(16#344C1#, 20), to_signed(16#344FB#, 20),
                                                                              to_signed(16#34535#, 20), to_signed(16#3456F#, 20), to_signed(16#345A9#, 20), to_signed(16#345E2#, 20),
                                                                              to_signed(16#3461C#, 20), to_signed(16#34656#, 20), to_signed(16#34690#, 20), to_signed(16#346C9#, 20),
                                                                              to_signed(16#34703#, 20), to_signed(16#3473D#, 20), to_signed(16#34776#, 20), to_signed(16#347B0#, 20),
                                                                              to_signed(16#347E9#, 20), to_signed(16#34823#, 20), to_signed(16#3485C#, 20), to_signed(16#34896#, 20),
                                                                              to_signed(16#348CF#, 20), to_signed(16#34908#, 20), to_signed(16#34942#, 20), to_signed(16#3497B#, 20),
                                                                              to_signed(16#349B4#, 20), to_signed(16#349EE#, 20), to_signed(16#34A27#, 20), to_signed(16#34A60#, 20),
                                                                              to_signed(16#34A99#, 20), to_signed(16#34AD2#, 20), to_signed(16#34B0B#, 20), to_signed(16#34B44#, 20),
                                                                              to_signed(16#34B7D#, 20), to_signed(16#34BB6#, 20), to_signed(16#34BEF#, 20), to_signed(16#34C28#, 20),
                                                                              to_signed(16#34C61#, 20), to_signed(16#34C9A#, 20), to_signed(16#34CD3#, 20), to_signed(16#34D0C#, 20),
                                                                              to_signed(16#34D44#, 20), to_signed(16#34D7D#, 20), to_signed(16#34DB6#, 20), to_signed(16#34DEE#, 20),
                                                                              to_signed(16#34E27#, 20), to_signed(16#34E60#, 20), to_signed(16#34E98#, 20), to_signed(16#34ED1#, 20),
                                                                              to_signed(16#34F09#, 20), to_signed(16#34F42#, 20), to_signed(16#34F7A#, 20), to_signed(16#34FB3#, 20),
                                                                              to_signed(16#34FEB#, 20), to_signed(16#35023#, 20), to_signed(16#3505C#, 20), to_signed(16#35094#, 20),
                                                                              to_signed(16#350CC#, 20), to_signed(16#35104#, 20), to_signed(16#3513D#, 20), to_signed(16#35175#, 20),
                                                                              to_signed(16#351AD#, 20), to_signed(16#351E5#, 20), to_signed(16#3521D#, 20), to_signed(16#35255#, 20),
                                                                              to_signed(16#3528D#, 20), to_signed(16#352C5#, 20), to_signed(16#352FD#, 20), to_signed(16#35335#, 20),
                                                                              to_signed(16#3536D#, 20), to_signed(16#353A5#, 20), to_signed(16#353DC#, 20), to_signed(16#35414#, 20),
                                                                              to_signed(16#3544C#, 20), to_signed(16#35484#, 20), to_signed(16#354BB#, 20), to_signed(16#354F3#, 20),
                                                                              to_signed(16#3552B#, 20), to_signed(16#35562#, 20), to_signed(16#3559A#, 20), to_signed(16#355D1#, 20),
                                                                              to_signed(16#35609#, 20), to_signed(16#35640#, 20), to_signed(16#35678#, 20), to_signed(16#356AF#, 20),
                                                                              to_signed(16#356E6#, 20), to_signed(16#3571E#, 20), to_signed(16#35755#, 20), to_signed(16#3578C#, 20),
                                                                              to_signed(16#357C3#, 20), to_signed(16#357FB#, 20), to_signed(16#35832#, 20), to_signed(16#35869#, 20),
                                                                              to_signed(16#358A0#, 20), to_signed(16#358D7#, 20), to_signed(16#3590E#, 20), to_signed(16#35945#, 20),
                                                                              to_signed(16#3597C#, 20), to_signed(16#359B3#, 20), to_signed(16#359EA#, 20), to_signed(16#35A21#, 20),
                                                                              to_signed(16#35A58#, 20), to_signed(16#35A8E#, 20), to_signed(16#35AC5#, 20), to_signed(16#35AFC#, 20),
                                                                              to_signed(16#35B33#, 20), to_signed(16#35B69#, 20), to_signed(16#35BA0#, 20), to_signed(16#35BD7#, 20),
                                                                              to_signed(16#35C0D#, 20), to_signed(16#35C44#, 20), to_signed(16#35C7A#, 20), to_signed(16#35CB1#, 20),
                                                                              to_signed(16#35CE7#, 20), to_signed(16#35D1E#, 20), to_signed(16#35D54#, 20), to_signed(16#35D8A#, 20),
                                                                              to_signed(16#35DC1#, 20), to_signed(16#35DF7#, 20), to_signed(16#35E2D#, 20), to_signed(16#35E63#, 20),
                                                                              to_signed(16#35E9A#, 20), to_signed(16#35ED0#, 20), to_signed(16#35F06#, 20), to_signed(16#35F3C#, 20),
                                                                              to_signed(16#35F72#, 20), to_signed(16#35FA8#, 20), to_signed(16#35FDE#, 20), to_signed(16#36014#, 20),
                                                                              to_signed(16#3604A#, 20), to_signed(16#36080#, 20), to_signed(16#360B6#, 20), to_signed(16#360EB#, 20),
                                                                              to_signed(16#36121#, 20), to_signed(16#36157#, 20), to_signed(16#3618D#, 20), to_signed(16#361C2#, 20),
                                                                              to_signed(16#361F8#, 20), to_signed(16#3622E#, 20), to_signed(16#36263#, 20), to_signed(16#36299#, 20),
                                                                              to_signed(16#362CF#, 20), to_signed(16#36304#, 20), to_signed(16#3633A#, 20), to_signed(16#3636F#, 20),
                                                                              to_signed(16#363A4#, 20), to_signed(16#363DA#, 20), to_signed(16#3640F#, 20), to_signed(16#36444#, 20),
                                                                              to_signed(16#3647A#, 20), to_signed(16#364AF#, 20), to_signed(16#364E4#, 20), to_signed(16#36519#, 20),
                                                                              to_signed(16#3654E#, 20), to_signed(16#36584#, 20), to_signed(16#365B9#, 20), to_signed(16#365EE#, 20),
                                                                              to_signed(16#36623#, 20), to_signed(16#36658#, 20), to_signed(16#3668D#, 20), to_signed(16#366C2#, 20),
                                                                              to_signed(16#366F6#, 20), to_signed(16#3672B#, 20), to_signed(16#36760#, 20), to_signed(16#36795#, 20),
                                                                              to_signed(16#367CA#, 20), to_signed(16#367FE#, 20), to_signed(16#36833#, 20), to_signed(16#36868#, 20),
                                                                              to_signed(16#3689C#, 20), to_signed(16#368D1#, 20), to_signed(16#36905#, 20), to_signed(16#3693A#, 20),
                                                                              to_signed(16#3696F#, 20), to_signed(16#369A3#, 20), to_signed(16#369D7#, 20), to_signed(16#36A0C#, 20),
                                                                              to_signed(16#36A40#, 20), to_signed(16#36A74#, 20), to_signed(16#36AA9#, 20), to_signed(16#36ADD#, 20),
                                                                              to_signed(16#36B11#, 20), to_signed(16#36B45#, 20), to_signed(16#36B7A#, 20), to_signed(16#36BAE#, 20),
                                                                              to_signed(16#36BE2#, 20), to_signed(16#36C16#, 20), to_signed(16#36C4A#, 20), to_signed(16#36C7E#, 20),
                                                                              to_signed(16#36CB2#, 20), to_signed(16#36CE6#, 20), to_signed(16#36D1A#, 20), to_signed(16#36D4E#, 20),
                                                                              to_signed(16#36D81#, 20), to_signed(16#36DB5#, 20), to_signed(16#36DE9#, 20), to_signed(16#36E1D#, 20),
                                                                              to_signed(16#36E50#, 20), to_signed(16#36E84#, 20), to_signed(16#36EB8#, 20), to_signed(16#36EEB#, 20),
                                                                              to_signed(16#36F1F#, 20), to_signed(16#36F52#, 20), to_signed(16#36F86#, 20), to_signed(16#36FB9#, 20),
                                                                              to_signed(16#36FED#, 20), to_signed(16#37020#, 20), to_signed(16#37054#, 20), to_signed(16#37087#, 20),
                                                                              to_signed(16#370BA#, 20), to_signed(16#370ED#, 20), to_signed(16#37121#, 20), to_signed(16#37154#, 20),
                                                                              to_signed(16#37187#, 20), to_signed(16#371BA#, 20), to_signed(16#371ED#, 20), to_signed(16#37220#, 20),
                                                                              to_signed(16#37253#, 20), to_signed(16#37286#, 20), to_signed(16#372B9#, 20), to_signed(16#372EC#, 20),
                                                                              to_signed(16#3731F#, 20), to_signed(16#37352#, 20), to_signed(16#37385#, 20), to_signed(16#373B8#, 20),
                                                                              to_signed(16#373EB#, 20), to_signed(16#3741D#, 20), to_signed(16#37450#, 20), to_signed(16#37483#, 20),
                                                                              to_signed(16#374B5#, 20), to_signed(16#374E8#, 20), to_signed(16#3751A#, 20), to_signed(16#3754D#, 20),
                                                                              to_signed(16#37580#, 20), to_signed(16#375B2#, 20), to_signed(16#375E4#, 20), to_signed(16#37617#, 20),
                                                                              to_signed(16#37649#, 20), to_signed(16#3767C#, 20), to_signed(16#376AE#, 20), to_signed(16#376E0#, 20),
                                                                              to_signed(16#37712#, 20), to_signed(16#37745#, 20), to_signed(16#37777#, 20), to_signed(16#377A9#, 20),
                                                                              to_signed(16#377DB#, 20), to_signed(16#3780D#, 20), to_signed(16#3783F#, 20), to_signed(16#37871#, 20),
                                                                              to_signed(16#378A3#, 20), to_signed(16#378D5#, 20), to_signed(16#37907#, 20), to_signed(16#37939#, 20),
                                                                              to_signed(16#3796B#, 20), to_signed(16#3799C#, 20), to_signed(16#379CE#, 20), to_signed(16#37A00#, 20),
                                                                              to_signed(16#37A32#, 20), to_signed(16#37A63#, 20), to_signed(16#37A95#, 20), to_signed(16#37AC7#, 20),
                                                                              to_signed(16#37AF8#, 20), to_signed(16#37B2A#, 20), to_signed(16#37B5B#, 20), to_signed(16#37B8D#, 20),
                                                                              to_signed(16#37BBE#, 20), to_signed(16#37BEF#, 20), to_signed(16#37C21#, 20), to_signed(16#37C52#, 20),
                                                                              to_signed(16#37C83#, 20), to_signed(16#37CB5#, 20), to_signed(16#37CE6#, 20), to_signed(16#37D17#, 20),
                                                                              to_signed(16#37D48#, 20), to_signed(16#37D79#, 20), to_signed(16#37DAB#, 20), to_signed(16#37DDC#, 20),
                                                                              to_signed(16#37E0D#, 20), to_signed(16#37E3E#, 20), to_signed(16#37E6F#, 20), to_signed(16#37EA0#, 20),
                                                                              to_signed(16#37ED0#, 20), to_signed(16#37F01#, 20), to_signed(16#37F32#, 20), to_signed(16#37F63#, 20),
                                                                              to_signed(16#37F94#, 20), to_signed(16#37FC4#, 20), to_signed(16#37FF5#, 20), to_signed(16#38026#, 20),
                                                                              to_signed(16#38056#, 20), to_signed(16#38087#, 20), to_signed(16#380B8#, 20), to_signed(16#380E8#, 20),
                                                                              to_signed(16#38119#, 20), to_signed(16#38149#, 20), to_signed(16#38179#, 20), to_signed(16#381AA#, 20),
                                                                              to_signed(16#381DA#, 20), to_signed(16#3820A#, 20), to_signed(16#3823B#, 20), to_signed(16#3826B#, 20),
                                                                              to_signed(16#3829B#, 20), to_signed(16#382CB#, 20), to_signed(16#382FC#, 20), to_signed(16#3832C#, 20),
                                                                              to_signed(16#3835C#, 20), to_signed(16#3838C#, 20), to_signed(16#383BC#, 20), to_signed(16#383EC#, 20),
                                                                              to_signed(16#3841C#, 20), to_signed(16#3844C#, 20), to_signed(16#3847C#, 20), to_signed(16#384AB#, 20),
                                                                              to_signed(16#384DB#, 20), to_signed(16#3850B#, 20), to_signed(16#3853B#, 20), to_signed(16#3856A#, 20),
                                                                              to_signed(16#3859A#, 20), to_signed(16#385CA#, 20), to_signed(16#385F9#, 20), to_signed(16#38629#, 20),
                                                                              to_signed(16#38659#, 20), to_signed(16#38688#, 20), to_signed(16#386B8#, 20), to_signed(16#386E7#, 20),
                                                                              to_signed(16#38716#, 20), to_signed(16#38746#, 20), to_signed(16#38775#, 20), to_signed(16#387A4#, 20),
                                                                              to_signed(16#387D4#, 20), to_signed(16#38803#, 20), to_signed(16#38832#, 20), to_signed(16#38861#, 20),
                                                                              to_signed(16#38890#, 20), to_signed(16#388BF#, 20), to_signed(16#388EF#, 20), to_signed(16#3891E#, 20),
                                                                              to_signed(16#3894D#, 20), to_signed(16#3897C#, 20), to_signed(16#389AA#, 20), to_signed(16#389D9#, 20),
                                                                              to_signed(16#38A08#, 20), to_signed(16#38A37#, 20), to_signed(16#38A66#, 20), to_signed(16#38A95#, 20),
                                                                              to_signed(16#38AC3#, 20), to_signed(16#38AF2#, 20), to_signed(16#38B21#, 20), to_signed(16#38B4F#, 20),
                                                                              to_signed(16#38B7E#, 20), to_signed(16#38BAC#, 20), to_signed(16#38BDB#, 20), to_signed(16#38C09#, 20),
                                                                              to_signed(16#38C38#, 20), to_signed(16#38C66#, 20), to_signed(16#38C95#, 20), to_signed(16#38CC3#, 20),
                                                                              to_signed(16#38CF1#, 20), to_signed(16#38D20#, 20), to_signed(16#38D4E#, 20), to_signed(16#38D7C#, 20),
                                                                              to_signed(16#38DAA#, 20), to_signed(16#38DD8#, 20), to_signed(16#38E07#, 20), to_signed(16#38E35#, 20),
                                                                              to_signed(16#38E63#, 20), to_signed(16#38E91#, 20), to_signed(16#38EBF#, 20), to_signed(16#38EED#, 20),
                                                                              to_signed(16#38F1B#, 20), to_signed(16#38F48#, 20), to_signed(16#38F76#, 20), to_signed(16#38FA4#, 20),
                                                                              to_signed(16#38FD2#, 20), to_signed(16#39000#, 20), to_signed(16#3902D#, 20), to_signed(16#3905B#, 20),
                                                                              to_signed(16#39089#, 20), to_signed(16#390B6#, 20), to_signed(16#390E4#, 20), to_signed(16#39111#, 20),
                                                                              to_signed(16#3913F#, 20), to_signed(16#3916C#, 20), to_signed(16#3919A#, 20), to_signed(16#391C7#, 20),
                                                                              to_signed(16#391F4#, 20), to_signed(16#39222#, 20), to_signed(16#3924F#, 20), to_signed(16#3927C#, 20),
                                                                              to_signed(16#392A9#, 20), to_signed(16#392D7#, 20), to_signed(16#39304#, 20), to_signed(16#39331#, 20),
                                                                              to_signed(16#3935E#, 20), to_signed(16#3938B#, 20), to_signed(16#393B8#, 20), to_signed(16#393E5#, 20),
                                                                              to_signed(16#39412#, 20), to_signed(16#3943F#, 20), to_signed(16#3946C#, 20), to_signed(16#39499#, 20),
                                                                              to_signed(16#394C5#, 20), to_signed(16#394F2#, 20), to_signed(16#3951F#, 20), to_signed(16#3954C#, 20),
                                                                              to_signed(16#39578#, 20), to_signed(16#395A5#, 20), to_signed(16#395D1#, 20), to_signed(16#395FE#, 20),
                                                                              to_signed(16#3962A#, 20), to_signed(16#39657#, 20), to_signed(16#39683#, 20), to_signed(16#396B0#, 20),
                                                                              to_signed(16#396DC#, 20), to_signed(16#39709#, 20), to_signed(16#39735#, 20), to_signed(16#39761#, 20),
                                                                              to_signed(16#3978D#, 20), to_signed(16#397BA#, 20), to_signed(16#397E6#, 20), to_signed(16#39812#, 20),
                                                                              to_signed(16#3983E#, 20), to_signed(16#3986A#, 20), to_signed(16#39896#, 20), to_signed(16#398C2#, 20),
                                                                              to_signed(16#398EE#, 20), to_signed(16#3991A#, 20), to_signed(16#39946#, 20), to_signed(16#39972#, 20),
                                                                              to_signed(16#3999E#, 20), to_signed(16#399CA#, 20), to_signed(16#399F5#, 20), to_signed(16#39A21#, 20),
                                                                              to_signed(16#39A4D#, 20), to_signed(16#39A78#, 20), to_signed(16#39AA4#, 20), to_signed(16#39AD0#, 20),
                                                                              to_signed(16#39AFB#, 20), to_signed(16#39B27#, 20), to_signed(16#39B52#, 20), to_signed(16#39B7E#, 20),
                                                                              to_signed(16#39BA9#, 20), to_signed(16#39BD4#, 20), to_signed(16#39C00#, 20), to_signed(16#39C2B#, 20),
                                                                              to_signed(16#39C56#, 20), to_signed(16#39C82#, 20), to_signed(16#39CAD#, 20), to_signed(16#39CD8#, 20),
                                                                              to_signed(16#39D03#, 20), to_signed(16#39D2E#, 20), to_signed(16#39D59#, 20), to_signed(16#39D84#, 20),
                                                                              to_signed(16#39DAF#, 20), to_signed(16#39DDA#, 20), to_signed(16#39E05#, 20), to_signed(16#39E30#, 20),
                                                                              to_signed(16#39E5B#, 20), to_signed(16#39E86#, 20), to_signed(16#39EB1#, 20), to_signed(16#39EDB#, 20),
                                                                              to_signed(16#39F06#, 20), to_signed(16#39F31#, 20), to_signed(16#39F5B#, 20), to_signed(16#39F86#, 20),
                                                                              to_signed(16#39FB1#, 20), to_signed(16#39FDB#, 20), to_signed(16#3A006#, 20), to_signed(16#3A030#, 20),
                                                                              to_signed(16#3A05B#, 20), to_signed(16#3A085#, 20), to_signed(16#3A0AF#, 20), to_signed(16#3A0DA#, 20),
                                                                              to_signed(16#3A104#, 20), to_signed(16#3A12E#, 20), to_signed(16#3A159#, 20), to_signed(16#3A183#, 20),
                                                                              to_signed(16#3A1AD#, 20), to_signed(16#3A1D7#, 20), to_signed(16#3A201#, 20), to_signed(16#3A22B#, 20),
                                                                              to_signed(16#3A255#, 20), to_signed(16#3A27F#, 20), to_signed(16#3A2A9#, 20), to_signed(16#3A2D3#, 20),
                                                                              to_signed(16#3A2FD#, 20), to_signed(16#3A327#, 20), to_signed(16#3A351#, 20), to_signed(16#3A37A#, 20),
                                                                              to_signed(16#3A3A4#, 20), to_signed(16#3A3CE#, 20), to_signed(16#3A3F7#, 20), to_signed(16#3A421#, 20),
                                                                              to_signed(16#3A44B#, 20), to_signed(16#3A474#, 20), to_signed(16#3A49E#, 20), to_signed(16#3A4C7#, 20),
                                                                              to_signed(16#3A4F1#, 20), to_signed(16#3A51A#, 20), to_signed(16#3A544#, 20), to_signed(16#3A56D#, 20),
                                                                              to_signed(16#3A596#, 20), to_signed(16#3A5C0#, 20), to_signed(16#3A5E9#, 20), to_signed(16#3A612#, 20),
                                                                              to_signed(16#3A63B#, 20), to_signed(16#3A664#, 20), to_signed(16#3A68D#, 20), to_signed(16#3A6B7#, 20),
                                                                              to_signed(16#3A6E0#, 20), to_signed(16#3A709#, 20), to_signed(16#3A732#, 20), to_signed(16#3A75A#, 20),
                                                                              to_signed(16#3A783#, 20), to_signed(16#3A7AC#, 20), to_signed(16#3A7D5#, 20), to_signed(16#3A7FE#, 20),
                                                                              to_signed(16#3A827#, 20), to_signed(16#3A84F#, 20), to_signed(16#3A878#, 20), to_signed(16#3A8A1#, 20),
                                                                              to_signed(16#3A8C9#, 20), to_signed(16#3A8F2#, 20), to_signed(16#3A91A#, 20), to_signed(16#3A943#, 20),
                                                                              to_signed(16#3A96B#, 20), to_signed(16#3A994#, 20), to_signed(16#3A9BC#, 20), to_signed(16#3A9E5#, 20),
                                                                              to_signed(16#3AA0D#, 20), to_signed(16#3AA35#, 20), to_signed(16#3AA5D#, 20), to_signed(16#3AA86#, 20),
                                                                              to_signed(16#3AAAE#, 20), to_signed(16#3AAD6#, 20), to_signed(16#3AAFE#, 20), to_signed(16#3AB26#, 20),
                                                                              to_signed(16#3AB4E#, 20), to_signed(16#3AB76#, 20), to_signed(16#3AB9E#, 20), to_signed(16#3ABC6#, 20),
                                                                              to_signed(16#3ABEE#, 20), to_signed(16#3AC16#, 20), to_signed(16#3AC3E#, 20), to_signed(16#3AC66#, 20),
                                                                              to_signed(16#3AC8D#, 20), to_signed(16#3ACB5#, 20), to_signed(16#3ACDD#, 20), to_signed(16#3AD05#, 20),
                                                                              to_signed(16#3AD2C#, 20), to_signed(16#3AD54#, 20), to_signed(16#3AD7B#, 20), to_signed(16#3ADA3#, 20),
                                                                              to_signed(16#3ADCA#, 20), to_signed(16#3ADF2#, 20), to_signed(16#3AE19#, 20), to_signed(16#3AE41#, 20),
                                                                              to_signed(16#3AE68#, 20), to_signed(16#3AE8F#, 20), to_signed(16#3AEB6#, 20), to_signed(16#3AEDE#, 20),
                                                                              to_signed(16#3AF05#, 20), to_signed(16#3AF2C#, 20), to_signed(16#3AF53#, 20), to_signed(16#3AF7A#, 20),
                                                                              to_signed(16#3AFA1#, 20), to_signed(16#3AFC8#, 20), to_signed(16#3AFEF#, 20), to_signed(16#3B016#, 20),
                                                                              to_signed(16#3B03D#, 20), to_signed(16#3B064#, 20), to_signed(16#3B08B#, 20), to_signed(16#3B0B2#, 20),
                                                                              to_signed(16#3B0D9#, 20), to_signed(16#3B0FF#, 20), to_signed(16#3B126#, 20), to_signed(16#3B14D#, 20),
                                                                              to_signed(16#3B173#, 20), to_signed(16#3B19A#, 20), to_signed(16#3B1C0#, 20), to_signed(16#3B1E7#, 20),
                                                                              to_signed(16#3B20D#, 20), to_signed(16#3B234#, 20), to_signed(16#3B25A#, 20), to_signed(16#3B281#, 20),
                                                                              to_signed(16#3B2A7#, 20), to_signed(16#3B2CD#, 20), to_signed(16#3B2F4#, 20), to_signed(16#3B31A#, 20),
                                                                              to_signed(16#3B340#, 20), to_signed(16#3B366#, 20), to_signed(16#3B38C#, 20), to_signed(16#3B3B3#, 20),
                                                                              to_signed(16#3B3D9#, 20), to_signed(16#3B3FF#, 20), to_signed(16#3B425#, 20), to_signed(16#3B44B#, 20),
                                                                              to_signed(16#3B470#, 20), to_signed(16#3B496#, 20), to_signed(16#3B4BC#, 20), to_signed(16#3B4E2#, 20),
                                                                              to_signed(16#3B508#, 20), to_signed(16#3B52E#, 20), to_signed(16#3B553#, 20), to_signed(16#3B579#, 20),
                                                                              to_signed(16#3B59F#, 20), to_signed(16#3B5C4#, 20), to_signed(16#3B5EA#, 20), to_signed(16#3B60F#, 20),
                                                                              to_signed(16#3B635#, 20), to_signed(16#3B65A#, 20), to_signed(16#3B680#, 20), to_signed(16#3B6A5#, 20),
                                                                              to_signed(16#3B6CA#, 20), to_signed(16#3B6F0#, 20), to_signed(16#3B715#, 20), to_signed(16#3B73A#, 20),
                                                                              to_signed(16#3B75F#, 20), to_signed(16#3B784#, 20), to_signed(16#3B7AA#, 20), to_signed(16#3B7CF#, 20),
                                                                              to_signed(16#3B7F4#, 20), to_signed(16#3B819#, 20), to_signed(16#3B83E#, 20), to_signed(16#3B863#, 20),
                                                                              to_signed(16#3B888#, 20), to_signed(16#3B8AD#, 20), to_signed(16#3B8D1#, 20), to_signed(16#3B8F6#, 20),
                                                                              to_signed(16#3B91B#, 20), to_signed(16#3B940#, 20), to_signed(16#3B964#, 20), to_signed(16#3B989#, 20),
                                                                              to_signed(16#3B9AE#, 20), to_signed(16#3B9D2#, 20), to_signed(16#3B9F7#, 20), to_signed(16#3BA1B#, 20),
                                                                              to_signed(16#3BA40#, 20), to_signed(16#3BA64#, 20), to_signed(16#3BA89#, 20), to_signed(16#3BAAD#, 20),
                                                                              to_signed(16#3BAD1#, 20), to_signed(16#3BAF6#, 20), to_signed(16#3BB1A#, 20), to_signed(16#3BB3E#, 20),
                                                                              to_signed(16#3BB62#, 20), to_signed(16#3BB87#, 20), to_signed(16#3BBAB#, 20), to_signed(16#3BBCF#, 20),
                                                                              to_signed(16#3BBF3#, 20), to_signed(16#3BC17#, 20), to_signed(16#3BC3B#, 20), to_signed(16#3BC5F#, 20),
                                                                              to_signed(16#3BC83#, 20), to_signed(16#3BCA7#, 20), to_signed(16#3BCCA#, 20), to_signed(16#3BCEE#, 20),
                                                                              to_signed(16#3BD12#, 20), to_signed(16#3BD36#, 20), to_signed(16#3BD59#, 20), to_signed(16#3BD7D#, 20),
                                                                              to_signed(16#3BDA1#, 20), to_signed(16#3BDC4#, 20), to_signed(16#3BDE8#, 20), to_signed(16#3BE0B#, 20),
                                                                              to_signed(16#3BE2F#, 20), to_signed(16#3BE52#, 20), to_signed(16#3BE76#, 20), to_signed(16#3BE99#, 20),
                                                                              to_signed(16#3BEBC#, 20), to_signed(16#3BEE0#, 20), to_signed(16#3BF03#, 20), to_signed(16#3BF26#, 20),
                                                                              to_signed(16#3BF49#, 20), to_signed(16#3BF6D#, 20), to_signed(16#3BF90#, 20), to_signed(16#3BFB3#, 20),
                                                                              to_signed(16#3BFD6#, 20), to_signed(16#3BFF9#, 20), to_signed(16#3C01C#, 20), to_signed(16#3C03F#, 20),
                                                                              to_signed(16#3C062#, 20), to_signed(16#3C084#, 20), to_signed(16#3C0A7#, 20), to_signed(16#3C0CA#, 20),
                                                                              to_signed(16#3C0ED#, 20), to_signed(16#3C110#, 20), to_signed(16#3C132#, 20), to_signed(16#3C155#, 20),
                                                                              to_signed(16#3C178#, 20), to_signed(16#3C19A#, 20), to_signed(16#3C1BD#, 20), to_signed(16#3C1DF#, 20),
                                                                              to_signed(16#3C202#, 20), to_signed(16#3C224#, 20), to_signed(16#3C246#, 20), to_signed(16#3C269#, 20),
                                                                              to_signed(16#3C28B#, 20), to_signed(16#3C2AD#, 20), to_signed(16#3C2D0#, 20), to_signed(16#3C2F2#, 20),
                                                                              to_signed(16#3C314#, 20), to_signed(16#3C336#, 20), to_signed(16#3C358#, 20), to_signed(16#3C37A#, 20),
                                                                              to_signed(16#3C39C#, 20), to_signed(16#3C3BE#, 20), to_signed(16#3C3E0#, 20), to_signed(16#3C402#, 20),
                                                                              to_signed(16#3C424#, 20), to_signed(16#3C446#, 20), to_signed(16#3C468#, 20), to_signed(16#3C48A#, 20),
                                                                              to_signed(16#3C4AB#, 20), to_signed(16#3C4CD#, 20), to_signed(16#3C4EF#, 20), to_signed(16#3C510#, 20),
                                                                              to_signed(16#3C532#, 20), to_signed(16#3C553#, 20), to_signed(16#3C575#, 20), to_signed(16#3C596#, 20),
                                                                              to_signed(16#3C5B8#, 20), to_signed(16#3C5D9#, 20), to_signed(16#3C5FB#, 20), to_signed(16#3C61C#, 20),
                                                                              to_signed(16#3C63D#, 20), to_signed(16#3C65F#, 20), to_signed(16#3C680#, 20), to_signed(16#3C6A1#, 20),
                                                                              to_signed(16#3C6C2#, 20), to_signed(16#3C6E3#, 20), to_signed(16#3C704#, 20), to_signed(16#3C725#, 20),
                                                                              to_signed(16#3C746#, 20), to_signed(16#3C767#, 20), to_signed(16#3C788#, 20), to_signed(16#3C7A9#, 20),
                                                                              to_signed(16#3C7CA#, 20), to_signed(16#3C7EB#, 20), to_signed(16#3C80C#, 20), to_signed(16#3C82D#, 20),
                                                                              to_signed(16#3C84D#, 20), to_signed(16#3C86E#, 20), to_signed(16#3C88F#, 20), to_signed(16#3C8AF#, 20),
                                                                              to_signed(16#3C8D0#, 20), to_signed(16#3C8F0#, 20), to_signed(16#3C911#, 20), to_signed(16#3C931#, 20),
                                                                              to_signed(16#3C952#, 20), to_signed(16#3C972#, 20), to_signed(16#3C993#, 20), to_signed(16#3C9B3#, 20),
                                                                              to_signed(16#3C9D3#, 20), to_signed(16#3C9F3#, 20), to_signed(16#3CA14#, 20), to_signed(16#3CA34#, 20),
                                                                              to_signed(16#3CA54#, 20), to_signed(16#3CA74#, 20), to_signed(16#3CA94#, 20), to_signed(16#3CAB4#, 20),
                                                                              to_signed(16#3CAD4#, 20), to_signed(16#3CAF4#, 20), to_signed(16#3CB14#, 20), to_signed(16#3CB34#, 20),
                                                                              to_signed(16#3CB54#, 20), to_signed(16#3CB73#, 20), to_signed(16#3CB93#, 20), to_signed(16#3CBB3#, 20),
                                                                              to_signed(16#3CBD3#, 20), to_signed(16#3CBF2#, 20), to_signed(16#3CC12#, 20), to_signed(16#3CC32#, 20),
                                                                              to_signed(16#3CC51#, 20), to_signed(16#3CC71#, 20), to_signed(16#3CC90#, 20), to_signed(16#3CCB0#, 20),
                                                                              to_signed(16#3CCCF#, 20), to_signed(16#3CCEE#, 20), to_signed(16#3CD0E#, 20), to_signed(16#3CD2D#, 20),
                                                                              to_signed(16#3CD4C#, 20), to_signed(16#3CD6B#, 20), to_signed(16#3CD8B#, 20), to_signed(16#3CDAA#, 20),
                                                                              to_signed(16#3CDC9#, 20), to_signed(16#3CDE8#, 20), to_signed(16#3CE07#, 20), to_signed(16#3CE26#, 20),
                                                                              to_signed(16#3CE45#, 20), to_signed(16#3CE64#, 20), to_signed(16#3CE83#, 20), to_signed(16#3CEA2#, 20),
                                                                              to_signed(16#3CEC0#, 20), to_signed(16#3CEDF#, 20), to_signed(16#3CEFE#, 20), to_signed(16#3CF1D#, 20),
                                                                              to_signed(16#3CF3B#, 20), to_signed(16#3CF5A#, 20), to_signed(16#3CF79#, 20), to_signed(16#3CF97#, 20),
                                                                              to_signed(16#3CFB6#, 20), to_signed(16#3CFD4#, 20), to_signed(16#3CFF3#, 20), to_signed(16#3D011#, 20),
                                                                              to_signed(16#3D02F#, 20), to_signed(16#3D04E#, 20), to_signed(16#3D06C#, 20), to_signed(16#3D08A#, 20),
                                                                              to_signed(16#3D0A9#, 20), to_signed(16#3D0C7#, 20), to_signed(16#3D0E5#, 20), to_signed(16#3D103#, 20),
                                                                              to_signed(16#3D121#, 20), to_signed(16#3D13F#, 20), to_signed(16#3D15D#, 20), to_signed(16#3D17B#, 20),
                                                                              to_signed(16#3D199#, 20), to_signed(16#3D1B7#, 20), to_signed(16#3D1D5#, 20), to_signed(16#3D1F3#, 20),
                                                                              to_signed(16#3D211#, 20), to_signed(16#3D22E#, 20), to_signed(16#3D24C#, 20), to_signed(16#3D26A#, 20),
                                                                              to_signed(16#3D287#, 20), to_signed(16#3D2A5#, 20), to_signed(16#3D2C2#, 20), to_signed(16#3D2E0#, 20),
                                                                              to_signed(16#3D2FE#, 20), to_signed(16#3D31B#, 20), to_signed(16#3D338#, 20), to_signed(16#3D356#, 20),
                                                                              to_signed(16#3D373#, 20), to_signed(16#3D390#, 20), to_signed(16#3D3AE#, 20), to_signed(16#3D3CB#, 20),
                                                                              to_signed(16#3D3E8#, 20), to_signed(16#3D405#, 20), to_signed(16#3D422#, 20), to_signed(16#3D440#, 20),
                                                                              to_signed(16#3D45D#, 20), to_signed(16#3D47A#, 20), to_signed(16#3D497#, 20), to_signed(16#3D4B4#, 20),
                                                                              to_signed(16#3D4D0#, 20), to_signed(16#3D4ED#, 20), to_signed(16#3D50A#, 20), to_signed(16#3D527#, 20),
                                                                              to_signed(16#3D544#, 20), to_signed(16#3D560#, 20), to_signed(16#3D57D#, 20), to_signed(16#3D59A#, 20),
                                                                              to_signed(16#3D5B6#, 20), to_signed(16#3D5D3#, 20), to_signed(16#3D5EF#, 20), to_signed(16#3D60C#, 20),
                                                                              to_signed(16#3D628#, 20), to_signed(16#3D645#, 20), to_signed(16#3D661#, 20), to_signed(16#3D67E#, 20),
                                                                              to_signed(16#3D69A#, 20), to_signed(16#3D6B6#, 20), to_signed(16#3D6D2#, 20), to_signed(16#3D6EF#, 20),
                                                                              to_signed(16#3D70B#, 20), to_signed(16#3D727#, 20), to_signed(16#3D743#, 20), to_signed(16#3D75F#, 20),
                                                                              to_signed(16#3D77B#, 20), to_signed(16#3D797#, 20), to_signed(16#3D7B3#, 20), to_signed(16#3D7CF#, 20),
                                                                              to_signed(16#3D7EB#, 20), to_signed(16#3D807#, 20), to_signed(16#3D822#, 20), to_signed(16#3D83E#, 20),
                                                                              to_signed(16#3D85A#, 20), to_signed(16#3D876#, 20), to_signed(16#3D891#, 20), to_signed(16#3D8AD#, 20),
                                                                              to_signed(16#3D8C8#, 20), to_signed(16#3D8E4#, 20), to_signed(16#3D8FF#, 20), to_signed(16#3D91B#, 20),
                                                                              to_signed(16#3D936#, 20), to_signed(16#3D952#, 20), to_signed(16#3D96D#, 20), to_signed(16#3D988#, 20),
                                                                              to_signed(16#3D9A4#, 20), to_signed(16#3D9BF#, 20), to_signed(16#3D9DA#, 20), to_signed(16#3D9F5#, 20),
                                                                              to_signed(16#3DA10#, 20), to_signed(16#3DA2C#, 20), to_signed(16#3DA47#, 20), to_signed(16#3DA62#, 20),
                                                                              to_signed(16#3DA7D#, 20), to_signed(16#3DA98#, 20), to_signed(16#3DAB2#, 20), to_signed(16#3DACD#, 20),
                                                                              to_signed(16#3DAE8#, 20), to_signed(16#3DB03#, 20), to_signed(16#3DB1E#, 20), to_signed(16#3DB38#, 20),
                                                                              to_signed(16#3DB53#, 20), to_signed(16#3DB6E#, 20), to_signed(16#3DB88#, 20), to_signed(16#3DBA3#, 20),
                                                                              to_signed(16#3DBBD#, 20), to_signed(16#3DBD8#, 20), to_signed(16#3DBF2#, 20), to_signed(16#3DC0D#, 20),
                                                                              to_signed(16#3DC27#, 20), to_signed(16#3DC42#, 20), to_signed(16#3DC5C#, 20), to_signed(16#3DC76#, 20),
                                                                              to_signed(16#3DC90#, 20), to_signed(16#3DCAB#, 20), to_signed(16#3DCC5#, 20), to_signed(16#3DCDF#, 20),
                                                                              to_signed(16#3DCF9#, 20), to_signed(16#3DD13#, 20), to_signed(16#3DD2D#, 20), to_signed(16#3DD47#, 20),
                                                                              to_signed(16#3DD61#, 20), to_signed(16#3DD7B#, 20), to_signed(16#3DD95#, 20), to_signed(16#3DDAF#, 20),
                                                                              to_signed(16#3DDC8#, 20), to_signed(16#3DDE2#, 20), to_signed(16#3DDFC#, 20), to_signed(16#3DE15#, 20),
                                                                              to_signed(16#3DE2F#, 20), to_signed(16#3DE49#, 20), to_signed(16#3DE62#, 20), to_signed(16#3DE7C#, 20),
                                                                              to_signed(16#3DE95#, 20), to_signed(16#3DEAF#, 20), to_signed(16#3DEC8#, 20), to_signed(16#3DEE2#, 20),
                                                                              to_signed(16#3DEFB#, 20), to_signed(16#3DF14#, 20), to_signed(16#3DF2D#, 20), to_signed(16#3DF47#, 20),
                                                                              to_signed(16#3DF60#, 20), to_signed(16#3DF79#, 20), to_signed(16#3DF92#, 20), to_signed(16#3DFAB#, 20),
                                                                              to_signed(16#3DFC4#, 20), to_signed(16#3DFDD#, 20), to_signed(16#3DFF6#, 20), to_signed(16#3E00F#, 20),
                                                                              to_signed(16#3E028#, 20), to_signed(16#3E041#, 20), to_signed(16#3E05A#, 20), to_signed(16#3E073#, 20),
                                                                              to_signed(16#3E08B#, 20), to_signed(16#3E0A4#, 20), to_signed(16#3E0BD#, 20), to_signed(16#3E0D5#, 20),
                                                                              to_signed(16#3E0EE#, 20), to_signed(16#3E106#, 20), to_signed(16#3E11F#, 20), to_signed(16#3E137#, 20),
                                                                              to_signed(16#3E150#, 20), to_signed(16#3E168#, 20), to_signed(16#3E181#, 20), to_signed(16#3E199#, 20),
                                                                              to_signed(16#3E1B1#, 20), to_signed(16#3E1CA#, 20), to_signed(16#3E1E2#, 20), to_signed(16#3E1FA#, 20),
                                                                              to_signed(16#3E212#, 20), to_signed(16#3E22A#, 20), to_signed(16#3E242#, 20), to_signed(16#3E25A#, 20),
                                                                              to_signed(16#3E272#, 20), to_signed(16#3E28A#, 20), to_signed(16#3E2A2#, 20), to_signed(16#3E2BA#, 20),
                                                                              to_signed(16#3E2D2#, 20), to_signed(16#3E2EA#, 20), to_signed(16#3E301#, 20), to_signed(16#3E319#, 20),
                                                                              to_signed(16#3E331#, 20), to_signed(16#3E349#, 20), to_signed(16#3E360#, 20), to_signed(16#3E378#, 20),
                                                                              to_signed(16#3E38F#, 20), to_signed(16#3E3A7#, 20), to_signed(16#3E3BE#, 20), to_signed(16#3E3D6#, 20),
                                                                              to_signed(16#3E3ED#, 20), to_signed(16#3E405#, 20), to_signed(16#3E41C#, 20), to_signed(16#3E433#, 20),
                                                                              to_signed(16#3E44A#, 20), to_signed(16#3E462#, 20), to_signed(16#3E479#, 20), to_signed(16#3E490#, 20),
                                                                              to_signed(16#3E4A7#, 20), to_signed(16#3E4BE#, 20), to_signed(16#3E4D5#, 20), to_signed(16#3E4EC#, 20),
                                                                              to_signed(16#3E503#, 20), to_signed(16#3E51A#, 20), to_signed(16#3E531#, 20), to_signed(16#3E548#, 20),
                                                                              to_signed(16#3E55E#, 20), to_signed(16#3E575#, 20), to_signed(16#3E58C#, 20), to_signed(16#3E5A3#, 20),
                                                                              to_signed(16#3E5B9#, 20), to_signed(16#3E5D0#, 20), to_signed(16#3E5E6#, 20), to_signed(16#3E5FD#, 20),
                                                                              to_signed(16#3E613#, 20), to_signed(16#3E62A#, 20), to_signed(16#3E640#, 20), to_signed(16#3E657#, 20),
                                                                              to_signed(16#3E66D#, 20), to_signed(16#3E683#, 20), to_signed(16#3E69A#, 20), to_signed(16#3E6B0#, 20),
                                                                              to_signed(16#3E6C6#, 20), to_signed(16#3E6DC#, 20), to_signed(16#3E6F2#, 20), to_signed(16#3E708#, 20),
                                                                              to_signed(16#3E71E#, 20), to_signed(16#3E734#, 20), to_signed(16#3E74A#, 20), to_signed(16#3E760#, 20),
                                                                              to_signed(16#3E776#, 20), to_signed(16#3E78C#, 20), to_signed(16#3E7A2#, 20), to_signed(16#3E7B8#, 20),
                                                                              to_signed(16#3E7CD#, 20), to_signed(16#3E7E3#, 20), to_signed(16#3E7F9#, 20), to_signed(16#3E80E#, 20),
                                                                              to_signed(16#3E824#, 20), to_signed(16#3E83A#, 20), to_signed(16#3E84F#, 20), to_signed(16#3E865#, 20),
                                                                              to_signed(16#3E87A#, 20), to_signed(16#3E88F#, 20), to_signed(16#3E8A5#, 20), to_signed(16#3E8BA#, 20),
                                                                              to_signed(16#3E8CF#, 20), to_signed(16#3E8E5#, 20), to_signed(16#3E8FA#, 20), to_signed(16#3E90F#, 20),
                                                                              to_signed(16#3E924#, 20), to_signed(16#3E939#, 20), to_signed(16#3E94E#, 20), to_signed(16#3E963#, 20),
                                                                              to_signed(16#3E978#, 20), to_signed(16#3E98D#, 20), to_signed(16#3E9A2#, 20), to_signed(16#3E9B7#, 20),
                                                                              to_signed(16#3E9CC#, 20), to_signed(16#3E9E1#, 20), to_signed(16#3E9F6#, 20), to_signed(16#3EA0A#, 20),
                                                                              to_signed(16#3EA1F#, 20), to_signed(16#3EA34#, 20), to_signed(16#3EA48#, 20), to_signed(16#3EA5D#, 20),
                                                                              to_signed(16#3EA71#, 20), to_signed(16#3EA86#, 20), to_signed(16#3EA9A#, 20), to_signed(16#3EAAF#, 20),
                                                                              to_signed(16#3EAC3#, 20), to_signed(16#3EAD8#, 20), to_signed(16#3EAEC#, 20), to_signed(16#3EB00#, 20),
                                                                              to_signed(16#3EB14#, 20), to_signed(16#3EB29#, 20), to_signed(16#3EB3D#, 20), to_signed(16#3EB51#, 20),
                                                                              to_signed(16#3EB65#, 20), to_signed(16#3EB79#, 20), to_signed(16#3EB8D#, 20), to_signed(16#3EBA1#, 20),
                                                                              to_signed(16#3EBB5#, 20), to_signed(16#3EBC9#, 20), to_signed(16#3EBDD#, 20), to_signed(16#3EBF0#, 20),
                                                                              to_signed(16#3EC04#, 20), to_signed(16#3EC18#, 20), to_signed(16#3EC2C#, 20), to_signed(16#3EC3F#, 20),
                                                                              to_signed(16#3EC53#, 20), to_signed(16#3EC67#, 20), to_signed(16#3EC7A#, 20), to_signed(16#3EC8E#, 20),
                                                                              to_signed(16#3ECA1#, 20), to_signed(16#3ECB5#, 20), to_signed(16#3ECC8#, 20), to_signed(16#3ECDB#, 20),
                                                                              to_signed(16#3ECEF#, 20), to_signed(16#3ED02#, 20), to_signed(16#3ED15#, 20), to_signed(16#3ED28#, 20),
                                                                              to_signed(16#3ED3C#, 20), to_signed(16#3ED4F#, 20), to_signed(16#3ED62#, 20), to_signed(16#3ED75#, 20),
                                                                              to_signed(16#3ED88#, 20), to_signed(16#3ED9B#, 20), to_signed(16#3EDAE#, 20), to_signed(16#3EDC1#, 20),
                                                                              to_signed(16#3EDD4#, 20), to_signed(16#3EDE6#, 20), to_signed(16#3EDF9#, 20), to_signed(16#3EE0C#, 20),
                                                                              to_signed(16#3EE1F#, 20), to_signed(16#3EE31#, 20), to_signed(16#3EE44#, 20), to_signed(16#3EE57#, 20),
                                                                              to_signed(16#3EE69#, 20), to_signed(16#3EE7C#, 20), to_signed(16#3EE8E#, 20), to_signed(16#3EEA1#, 20),
                                                                              to_signed(16#3EEB3#, 20), to_signed(16#3EEC6#, 20), to_signed(16#3EED8#, 20), to_signed(16#3EEEA#, 20),
                                                                              to_signed(16#3EEFD#, 20), to_signed(16#3EF0F#, 20), to_signed(16#3EF21#, 20), to_signed(16#3EF33#, 20),
                                                                              to_signed(16#3EF45#, 20), to_signed(16#3EF57#, 20), to_signed(16#3EF69#, 20), to_signed(16#3EF7B#, 20),
                                                                              to_signed(16#3EF8D#, 20), to_signed(16#3EF9F#, 20), to_signed(16#3EFB1#, 20), to_signed(16#3EFC3#, 20),
                                                                              to_signed(16#3EFD5#, 20), to_signed(16#3EFE7#, 20), to_signed(16#3EFF8#, 20), to_signed(16#3F00A#, 20),
                                                                              to_signed(16#3F01C#, 20), to_signed(16#3F02D#, 20), to_signed(16#3F03F#, 20), to_signed(16#3F050#, 20),
                                                                              to_signed(16#3F062#, 20), to_signed(16#3F073#, 20), to_signed(16#3F085#, 20), to_signed(16#3F096#, 20),
                                                                              to_signed(16#3F0A8#, 20), to_signed(16#3F0B9#, 20), to_signed(16#3F0CA#, 20), to_signed(16#3F0DB#, 20),
                                                                              to_signed(16#3F0ED#, 20), to_signed(16#3F0FE#, 20), to_signed(16#3F10F#, 20), to_signed(16#3F120#, 20),
                                                                              to_signed(16#3F131#, 20), to_signed(16#3F142#, 20), to_signed(16#3F153#, 20), to_signed(16#3F164#, 20),
                                                                              to_signed(16#3F175#, 20), to_signed(16#3F186#, 20), to_signed(16#3F197#, 20), to_signed(16#3F1A7#, 20),
                                                                              to_signed(16#3F1B8#, 20), to_signed(16#3F1C9#, 20), to_signed(16#3F1DA#, 20), to_signed(16#3F1EA#, 20),
                                                                              to_signed(16#3F1FB#, 20), to_signed(16#3F20B#, 20), to_signed(16#3F21C#, 20), to_signed(16#3F22C#, 20),
                                                                              to_signed(16#3F23D#, 20), to_signed(16#3F24D#, 20), to_signed(16#3F25E#, 20), to_signed(16#3F26E#, 20),
                                                                              to_signed(16#3F27E#, 20), to_signed(16#3F28E#, 20), to_signed(16#3F29F#, 20), to_signed(16#3F2AF#, 20),
                                                                              to_signed(16#3F2BF#, 20), to_signed(16#3F2CF#, 20), to_signed(16#3F2DF#, 20), to_signed(16#3F2EF#, 20),
                                                                              to_signed(16#3F2FF#, 20), to_signed(16#3F30F#, 20), to_signed(16#3F31F#, 20), to_signed(16#3F32F#, 20),
                                                                              to_signed(16#3F33F#, 20), to_signed(16#3F34F#, 20), to_signed(16#3F35E#, 20), to_signed(16#3F36E#, 20),
                                                                              to_signed(16#3F37E#, 20), to_signed(16#3F38D#, 20), to_signed(16#3F39D#, 20), to_signed(16#3F3AD#, 20),
                                                                              to_signed(16#3F3BC#, 20), to_signed(16#3F3CC#, 20), to_signed(16#3F3DB#, 20), to_signed(16#3F3EA#, 20),
                                                                              to_signed(16#3F3FA#, 20), to_signed(16#3F409#, 20), to_signed(16#3F418#, 20), to_signed(16#3F428#, 20),
                                                                              to_signed(16#3F437#, 20), to_signed(16#3F446#, 20), to_signed(16#3F455#, 20), to_signed(16#3F464#, 20),
                                                                              to_signed(16#3F473#, 20), to_signed(16#3F482#, 20), to_signed(16#3F491#, 20), to_signed(16#3F4A0#, 20),
                                                                              to_signed(16#3F4AF#, 20), to_signed(16#3F4BE#, 20), to_signed(16#3F4CD#, 20), to_signed(16#3F4DC#, 20),
                                                                              to_signed(16#3F4EB#, 20), to_signed(16#3F4F9#, 20), to_signed(16#3F508#, 20), to_signed(16#3F517#, 20),
                                                                              to_signed(16#3F525#, 20), to_signed(16#3F534#, 20), to_signed(16#3F543#, 20), to_signed(16#3F551#, 20),
                                                                              to_signed(16#3F55F#, 20), to_signed(16#3F56E#, 20), to_signed(16#3F57C#, 20), to_signed(16#3F58B#, 20),
                                                                              to_signed(16#3F599#, 20), to_signed(16#3F5A7#, 20), to_signed(16#3F5B5#, 20), to_signed(16#3F5C4#, 20),
                                                                              to_signed(16#3F5D2#, 20), to_signed(16#3F5E0#, 20), to_signed(16#3F5EE#, 20), to_signed(16#3F5FC#, 20),
                                                                              to_signed(16#3F60A#, 20), to_signed(16#3F618#, 20), to_signed(16#3F626#, 20), to_signed(16#3F634#, 20),
                                                                              to_signed(16#3F642#, 20), to_signed(16#3F650#, 20), to_signed(16#3F65D#, 20), to_signed(16#3F66B#, 20),
                                                                              to_signed(16#3F679#, 20), to_signed(16#3F686#, 20), to_signed(16#3F694#, 20), to_signed(16#3F6A2#, 20),
                                                                              to_signed(16#3F6AF#, 20), to_signed(16#3F6BD#, 20), to_signed(16#3F6CA#, 20), to_signed(16#3F6D8#, 20),
                                                                              to_signed(16#3F6E5#, 20), to_signed(16#3F6F2#, 20), to_signed(16#3F700#, 20), to_signed(16#3F70D#, 20),
                                                                              to_signed(16#3F71A#, 20), to_signed(16#3F727#, 20), to_signed(16#3F735#, 20), to_signed(16#3F742#, 20),
                                                                              to_signed(16#3F74F#, 20), to_signed(16#3F75C#, 20), to_signed(16#3F769#, 20), to_signed(16#3F776#, 20),
                                                                              to_signed(16#3F783#, 20), to_signed(16#3F790#, 20), to_signed(16#3F79D#, 20), to_signed(16#3F7A9#, 20),
                                                                              to_signed(16#3F7B6#, 20), to_signed(16#3F7C3#, 20), to_signed(16#3F7D0#, 20), to_signed(16#3F7DC#, 20),
                                                                              to_signed(16#3F7E9#, 20), to_signed(16#3F7F5#, 20), to_signed(16#3F802#, 20), to_signed(16#3F80F#, 20),
                                                                              to_signed(16#3F81B#, 20), to_signed(16#3F827#, 20), to_signed(16#3F834#, 20), to_signed(16#3F840#, 20),
                                                                              to_signed(16#3F84D#, 20), to_signed(16#3F859#, 20), to_signed(16#3F865#, 20), to_signed(16#3F871#, 20),
                                                                              to_signed(16#3F87D#, 20), to_signed(16#3F88A#, 20), to_signed(16#3F896#, 20), to_signed(16#3F8A2#, 20),
                                                                              to_signed(16#3F8AE#, 20), to_signed(16#3F8BA#, 20), to_signed(16#3F8C6#, 20), to_signed(16#3F8D2#, 20),
                                                                              to_signed(16#3F8DD#, 20), to_signed(16#3F8E9#, 20), to_signed(16#3F8F5#, 20), to_signed(16#3F901#, 20),
                                                                              to_signed(16#3F90D#, 20), to_signed(16#3F918#, 20), to_signed(16#3F924#, 20), to_signed(16#3F92F#, 20),
                                                                              to_signed(16#3F93B#, 20), to_signed(16#3F947#, 20), to_signed(16#3F952#, 20), to_signed(16#3F95D#, 20),
                                                                              to_signed(16#3F969#, 20), to_signed(16#3F974#, 20), to_signed(16#3F980#, 20), to_signed(16#3F98B#, 20),
                                                                              to_signed(16#3F996#, 20), to_signed(16#3F9A1#, 20), to_signed(16#3F9AD#, 20), to_signed(16#3F9B8#, 20),
                                                                              to_signed(16#3F9C3#, 20), to_signed(16#3F9CE#, 20), to_signed(16#3F9D9#, 20), to_signed(16#3F9E4#, 20),
                                                                              to_signed(16#3F9EF#, 20), to_signed(16#3F9FA#, 20), to_signed(16#3FA05#, 20), to_signed(16#3FA0F#, 20),
                                                                              to_signed(16#3FA1A#, 20), to_signed(16#3FA25#, 20), to_signed(16#3FA30#, 20), to_signed(16#3FA3A#, 20),
                                                                              to_signed(16#3FA45#, 20), to_signed(16#3FA50#, 20), to_signed(16#3FA5A#, 20), to_signed(16#3FA65#, 20),
                                                                              to_signed(16#3FA6F#, 20), to_signed(16#3FA7A#, 20), to_signed(16#3FA84#, 20), to_signed(16#3FA8E#, 20),
                                                                              to_signed(16#3FA99#, 20), to_signed(16#3FAA3#, 20), to_signed(16#3FAAD#, 20), to_signed(16#3FAB7#, 20),
                                                                              to_signed(16#3FAC2#, 20), to_signed(16#3FACC#, 20), to_signed(16#3FAD6#, 20), to_signed(16#3FAE0#, 20),
                                                                              to_signed(16#3FAEA#, 20), to_signed(16#3FAF4#, 20), to_signed(16#3FAFE#, 20), to_signed(16#3FB08#, 20),
                                                                              to_signed(16#3FB12#, 20), to_signed(16#3FB1C#, 20), to_signed(16#3FB25#, 20), to_signed(16#3FB2F#, 20),
                                                                              to_signed(16#3FB39#, 20), to_signed(16#3FB42#, 20), to_signed(16#3FB4C#, 20), to_signed(16#3FB56#, 20),
                                                                              to_signed(16#3FB5F#, 20), to_signed(16#3FB69#, 20), to_signed(16#3FB72#, 20), to_signed(16#3FB7C#, 20),
                                                                              to_signed(16#3FB85#, 20), to_signed(16#3FB8F#, 20), to_signed(16#3FB98#, 20), to_signed(16#3FBA1#, 20),
                                                                              to_signed(16#3FBAA#, 20), to_signed(16#3FBB4#, 20), to_signed(16#3FBBD#, 20), to_signed(16#3FBC6#, 20),
                                                                              to_signed(16#3FBCF#, 20), to_signed(16#3FBD8#, 20), to_signed(16#3FBE1#, 20), to_signed(16#3FBEA#, 20),
                                                                              to_signed(16#3FBF3#, 20), to_signed(16#3FBFC#, 20), to_signed(16#3FC05#, 20), to_signed(16#3FC0E#, 20),
                                                                              to_signed(16#3FC17#, 20), to_signed(16#3FC1F#, 20), to_signed(16#3FC28#, 20), to_signed(16#3FC31#, 20),
                                                                              to_signed(16#3FC39#, 20), to_signed(16#3FC42#, 20), to_signed(16#3FC4B#, 20), to_signed(16#3FC53#, 20),
                                                                              to_signed(16#3FC5C#, 20), to_signed(16#3FC64#, 20), to_signed(16#3FC6C#, 20), to_signed(16#3FC75#, 20),
                                                                              to_signed(16#3FC7D#, 20), to_signed(16#3FC85#, 20), to_signed(16#3FC8E#, 20), to_signed(16#3FC96#, 20),
                                                                              to_signed(16#3FC9E#, 20), to_signed(16#3FCA6#, 20), to_signed(16#3FCAE#, 20), to_signed(16#3FCB6#, 20),
                                                                              to_signed(16#3FCBE#, 20), to_signed(16#3FCC6#, 20), to_signed(16#3FCCE#, 20), to_signed(16#3FCD6#, 20),
                                                                              to_signed(16#3FCDE#, 20), to_signed(16#3FCE6#, 20), to_signed(16#3FCEE#, 20), to_signed(16#3FCF6#, 20),
                                                                              to_signed(16#3FCFD#, 20), to_signed(16#3FD05#, 20), to_signed(16#3FD0D#, 20), to_signed(16#3FD14#, 20),
                                                                              to_signed(16#3FD1C#, 20), to_signed(16#3FD23#, 20), to_signed(16#3FD2B#, 20), to_signed(16#3FD32#, 20),
                                                                              to_signed(16#3FD3A#, 20), to_signed(16#3FD41#, 20), to_signed(16#3FD48#, 20), to_signed(16#3FD50#, 20),
                                                                              to_signed(16#3FD57#, 20), to_signed(16#3FD5E#, 20), to_signed(16#3FD65#, 20), to_signed(16#3FD6D#, 20),
                                                                              to_signed(16#3FD74#, 20), to_signed(16#3FD7B#, 20), to_signed(16#3FD82#, 20), to_signed(16#3FD89#, 20),
                                                                              to_signed(16#3FD90#, 20), to_signed(16#3FD97#, 20), to_signed(16#3FD9D#, 20), to_signed(16#3FDA4#, 20),
                                                                              to_signed(16#3FDAB#, 20), to_signed(16#3FDB2#, 20), to_signed(16#3FDB9#, 20), to_signed(16#3FDBF#, 20),
                                                                              to_signed(16#3FDC6#, 20), to_signed(16#3FDCD#, 20), to_signed(16#3FDD3#, 20), to_signed(16#3FDDA#, 20),
                                                                              to_signed(16#3FDE0#, 20), to_signed(16#3FDE7#, 20), to_signed(16#3FDED#, 20), to_signed(16#3FDF3#, 20),
                                                                              to_signed(16#3FDFA#, 20), to_signed(16#3FE00#, 20), to_signed(16#3FE06#, 20), to_signed(16#3FE0C#, 20),
                                                                              to_signed(16#3FE13#, 20), to_signed(16#3FE19#, 20), to_signed(16#3FE1F#, 20), to_signed(16#3FE25#, 20),
                                                                              to_signed(16#3FE2B#, 20), to_signed(16#3FE31#, 20), to_signed(16#3FE37#, 20), to_signed(16#3FE3D#, 20),
                                                                              to_signed(16#3FE43#, 20), to_signed(16#3FE49#, 20), to_signed(16#3FE4E#, 20), to_signed(16#3FE54#, 20),
                                                                              to_signed(16#3FE5A#, 20), to_signed(16#3FE60#, 20), to_signed(16#3FE65#, 20), to_signed(16#3FE6B#, 20),
                                                                              to_signed(16#3FE70#, 20), to_signed(16#3FE76#, 20), to_signed(16#3FE7B#, 20), to_signed(16#3FE81#, 20),
                                                                              to_signed(16#3FE86#, 20), to_signed(16#3FE8C#, 20), to_signed(16#3FE91#, 20), to_signed(16#3FE96#, 20),
                                                                              to_signed(16#3FE9C#, 20), to_signed(16#3FEA1#, 20), to_signed(16#3FEA6#, 20), to_signed(16#3FEAB#, 20),
                                                                              to_signed(16#3FEB0#, 20), to_signed(16#3FEB5#, 20), to_signed(16#3FEBA#, 20), to_signed(16#3FEBF#, 20),
                                                                              to_signed(16#3FEC4#, 20), to_signed(16#3FEC9#, 20), to_signed(16#3FECE#, 20), to_signed(16#3FED3#, 20),
                                                                              to_signed(16#3FED8#, 20), to_signed(16#3FEDC#, 20), to_signed(16#3FEE1#, 20), to_signed(16#3FEE6#, 20),
                                                                              to_signed(16#3FEEA#, 20), to_signed(16#3FEEF#, 20), to_signed(16#3FEF4#, 20), to_signed(16#3FEF8#, 20),
                                                                              to_signed(16#3FEFD#, 20), to_signed(16#3FF01#, 20), to_signed(16#3FF06#, 20), to_signed(16#3FF0A#, 20),
                                                                              to_signed(16#3FF0E#, 20), to_signed(16#3FF13#, 20), to_signed(16#3FF17#, 20), to_signed(16#3FF1B#, 20),
                                                                              to_signed(16#3FF1F#, 20), to_signed(16#3FF23#, 20), to_signed(16#3FF27#, 20), to_signed(16#3FF2C#, 20),
                                                                              to_signed(16#3FF30#, 20), to_signed(16#3FF34#, 20), to_signed(16#3FF37#, 20), to_signed(16#3FF3B#, 20),
                                                                              to_signed(16#3FF3F#, 20), to_signed(16#3FF43#, 20), to_signed(16#3FF47#, 20), to_signed(16#3FF4B#, 20),
                                                                              to_signed(16#3FF4E#, 20), to_signed(16#3FF52#, 20), to_signed(16#3FF56#, 20), to_signed(16#3FF59#, 20),
                                                                              to_signed(16#3FF5D#, 20), to_signed(16#3FF60#, 20), to_signed(16#3FF64#, 20), to_signed(16#3FF67#, 20),
                                                                              to_signed(16#3FF6B#, 20), to_signed(16#3FF6E#, 20), to_signed(16#3FF71#, 20), to_signed(16#3FF75#, 20),
                                                                              to_signed(16#3FF78#, 20), to_signed(16#3FF7B#, 20), to_signed(16#3FF7E#, 20), to_signed(16#3FF82#, 20),
                                                                              to_signed(16#3FF85#, 20), to_signed(16#3FF88#, 20), to_signed(16#3FF8B#, 20), to_signed(16#3FF8E#, 20),
                                                                              to_signed(16#3FF91#, 20), to_signed(16#3FF94#, 20), to_signed(16#3FF96#, 20), to_signed(16#3FF99#, 20),
                                                                              to_signed(16#3FF9C#, 20), to_signed(16#3FF9F#, 20), to_signed(16#3FFA2#, 20), to_signed(16#3FFA4#, 20),
                                                                              to_signed(16#3FFA7#, 20), to_signed(16#3FFA9#, 20), to_signed(16#3FFAC#, 20), to_signed(16#3FFAF#, 20),
                                                                              to_signed(16#3FFB1#, 20), to_signed(16#3FFB3#, 20), to_signed(16#3FFB6#, 20), to_signed(16#3FFB8#, 20),
                                                                              to_signed(16#3FFBB#, 20), to_signed(16#3FFBD#, 20), to_signed(16#3FFBF#, 20), to_signed(16#3FFC1#, 20),
                                                                              to_signed(16#3FFC4#, 20), to_signed(16#3FFC6#, 20), to_signed(16#3FFC8#, 20), to_signed(16#3FFCA#, 20),
                                                                              to_signed(16#3FFCC#, 20), to_signed(16#3FFCE#, 20), to_signed(16#3FFD0#, 20), to_signed(16#3FFD2#, 20),
                                                                              to_signed(16#3FFD4#, 20), to_signed(16#3FFD5#, 20), to_signed(16#3FFD7#, 20), to_signed(16#3FFD9#, 20),
                                                                              to_signed(16#3FFDB#, 20), to_signed(16#3FFDC#, 20), to_signed(16#3FFDE#, 20), to_signed(16#3FFE0#, 20),
                                                                              to_signed(16#3FFE1#, 20), to_signed(16#3FFE3#, 20), to_signed(16#3FFE4#, 20), to_signed(16#3FFE6#, 20),
                                                                              to_signed(16#3FFE7#, 20), to_signed(16#3FFE8#, 20), to_signed(16#3FFEA#, 20), to_signed(16#3FFEB#, 20),
                                                                              to_signed(16#3FFEC#, 20), to_signed(16#3FFED#, 20), to_signed(16#3FFEF#, 20), to_signed(16#3FFF0#, 20),
                                                                              to_signed(16#3FFF1#, 20), to_signed(16#3FFF2#, 20), to_signed(16#3FFF3#, 20), to_signed(16#3FFF4#, 20),
                                                                              to_signed(16#3FFF5#, 20), to_signed(16#3FFF6#, 20), to_signed(16#3FFF7#, 20), to_signed(16#3FFF7#, 20),
                                                                              to_signed(16#3FFF8#, 20), to_signed(16#3FFF9#, 20), to_signed(16#3FFFA#, 20), to_signed(16#3FFFA#, 20),
                                                                              to_signed(16#3FFFB#, 20), to_signed(16#3FFFC#, 20), to_signed(16#3FFFC#, 20), to_signed(16#3FFFD#, 20),
                                                                              to_signed(16#3FFFD#, 20), to_signed(16#3FFFE#, 20), to_signed(16#3FFFE#, 20), to_signed(16#3FFFE#, 20),
                                                                              to_signed(16#3FFFF#, 20), to_signed(16#3FFFF#, 20), to_signed(16#3FFFF#, 20), to_signed(16#40000#, 20),
                                                                              to_signed(16#40000#, 20), to_signed(16#40000#, 20), to_signed(16#40000#, 20), to_signed(16#40000#, 20) );  -- sfix20 [4096]
  CONSTANT table_data_2                   : vector_of_unsigned5(0 TO 4095) := ( to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#01000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00111#, 5), to_unsigned(2#00111#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00110#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5), to_unsigned(2#00101#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00100#, 5), to_unsigned(2#00100#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5), to_unsigned(2#00011#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00010#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5), to_unsigned(2#00001#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5),
                                                                               to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5), to_unsigned(2#00000#, 5) );  -- ufix5 [4096]

  -- Signals
  SIGNAL lutaddr_unsigned                 : unsigned(17 DOWNTO 0);  -- ufix18
  SIGNAL lutaddrInReg                     : unsigned(17 DOWNTO 0);  -- ufix18
  SIGNAL lut1addr                         : unsigned(11 DOWNTO 0);  -- ufix12
  SIGNAL Lookup_Table1_k                  : unsigned(11 DOWNTO 0);  -- ufix12
  SIGNAL lut1out                          : signed(19 DOWNTO 0);  -- sfix20_En18
  SIGNAL lut1out_rstnonereg               : signed(19 DOWNTO 0);  -- sfix20_En18
  SIGNAL lut2addrp1                       : unsigned(5 DOWNTO 0);  -- ufix6
  SIGNAL lut2addrp2                       : unsigned(5 DOWNTO 0);  -- ufix6
  SIGNAL lut2addr                         : unsigned(11 DOWNTO 0);  -- ufix12
  SIGNAL Lookup_Table2_k                  : unsigned(11 DOWNTO 0);  -- ufix12
  SIGNAL lut2out                          : unsigned(4 DOWNTO 0);  -- ufix5_En5
  SIGNAL lut2out_rstnonereg               : unsigned(4 DOWNTO 0);  -- ufix5_En5
  SIGNAL lut1outreg                       : signed(19 DOWNTO 0);  -- sfix20_En18
  SIGNAL lut2outreg                       : unsigned(4 DOWNTO 0);  -- ufix5_En5
  SIGNAL lut2out_extend                   : signed(19 DOWNTO 0);  -- sfix20_En18
  SIGNAL lut2out_sf                       : signed(19 DOWNTO 0);  -- sfix20_En18
  SIGNAL adder_add_cast                   : signed(20 DOWNTO 0);  -- sfix21_En18
  SIGNAL adder_add_cast_1                 : signed(20 DOWNTO 0);  -- sfix21_En18
  SIGNAL adder_add_temp                   : signed(20 DOWNTO 0);  -- sfix21_En18
  SIGNAL addlutouts                       : signed(19 DOWNTO 0);  -- sfix20_En18
  SIGNAL lutoutput_tmp                    : signed(19 DOWNTO 0);  -- sfix20_En18

BEGIN
  lutaddr_unsigned <= unsigned(lutaddr);

  -- Look up table address input register
  LUTaddrRegister_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        lutaddrInReg <= to_unsigned(2#000000000000000000#, 18);
      ELSIF enb = '1' THEN
        lutaddrInReg <= lutaddr_unsigned;
      END IF;
    END IF;
  END PROCESS LUTaddrRegister_process;


  -- Lookup table 1 address
  lut1addr <= lutaddrInReg(17 DOWNTO 6);

  -- Quarter sine wave table-Part1
  
  Lookup_Table1_k <= to_unsigned(2#000000000000#, 12) WHEN lut1addr <= 0 ELSE
      to_unsigned(2#111111111111#, 12) WHEN lut1addr >= 4095 ELSE
      lut1addr;
  lut1out <= table_data(to_integer(Lookup_Table1_k));

  -- Look up table1 output register-ResetNone
  LUT1outRegister_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
        lut1out_rstnonereg <= lut1out;
      END IF;
    END IF;
  END PROCESS LUT1outRegister_process;


  lut2addrp1 <= lutaddrInReg(17 DOWNTO 12);

  lut2addrp2 <= lutaddrInReg(5 DOWNTO 0);

  -- Lookup table 2 address
  lut2addr <= lut2addrp1 & lut2addrp2;

  -- Quarter Sine Wave Table-Part2
  
  Lookup_Table2_k <= to_unsigned(2#000000000000#, 12) WHEN lut2addr <= 0 ELSE
      to_unsigned(2#111111111111#, 12) WHEN lut2addr >= 4095 ELSE
      lut2addr;
  lut2out <= table_data_2(to_integer(Lookup_Table2_k));

  -- Look up table2 output register-ResetNone
  LUT2outRegister_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
        lut2out_rstnonereg <= lut2out;
      END IF;
    END IF;
  END PROCESS LUT2outRegister_process;


  LUToutRegister_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        lut1outreg <= to_signed(16#00000#, 20);
      ELSIF enb = '1' THEN
        lut1outreg <= lut1out_rstnonereg;
      END IF;
    END IF;
  END PROCESS LUToutRegister_process;


  LUToutRegister_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        lut2outreg <= to_unsigned(2#00000#, 5);
      ELSIF enb = '1' THEN
        lut2outreg <= lut2out_rstnonereg;
      END IF;
    END IF;
  END PROCESS LUToutRegister_1_process;


  lut2out_extend <= signed(resize(lut2outreg & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0', 20));

  -- Shift look up table 2 outputs
  lut2out_sf <= lut2out_extend srl 10;

  -- Compute look up table output
  adder_add_cast <= resize(lut1outreg, 21);
  adder_add_cast_1 <= resize(lut2out_sf, 21);
  adder_add_temp <= adder_add_cast + adder_add_cast_1;
  
  addlutouts <= X"7FFFF" WHEN (adder_add_temp(20) = '0') AND (adder_add_temp(19) /= '0') ELSE
      X"80000" WHEN (adder_add_temp(20) = '1') AND (adder_add_temp(19) /= '1') ELSE
      adder_add_temp(19 DOWNTO 0);

  -- Look up table output register
  LUToutRegister_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        lutoutput_tmp <= to_signed(16#00000#, 20);
      ELSIF enb = '1' THEN
        lutoutput_tmp <= addlutouts;
      END IF;
    END IF;
  END PROCESS LUToutRegister_2_process;


  lutoutput <= std_logic_vector(lutoutput_tmp);

END rtl;

